-- DVBT2_mod.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DVBT2_mod is
	port (
		baseband_i       : out std_logic_vector(13 downto 0);                    --      Baseband.i
		baseband_q       : out std_logic_vector(13 downto 0);                    --              .q
		baseband_valid   : out std_logic;                                        --              .valid
		fft_wr_addr      : out std_logic_vector(18 downto 0);                    --           QDR.fft_wr_addr
		fft_wr_data      : out std_logic_vector(35 downto 0);                    --              .fft_wr_data
		fft_wr_ena       : out std_logic;                                        --              .fft_wr_ena
		fft_rd_addr      : out std_logic_vector(18 downto 0);                    --              .fft_rd_addr
		fft_rd_data      : in  std_logic_vector(35 downto 0) := (others => '0'); --              .fft_rd_data
		osg_wr_addr      : out std_logic_vector(18 downto 0);                    --              .osg_wr_addr
		osg_wr_data      : out std_logic_vector(35 downto 0);                    --              .osg_wr_data
		osg_wr_ena       : out std_logic;                                        --              .osg_wr_ena
		osg_rd_addr      : out std_logic_vector(18 downto 0);                    --              .osg_rd_addr
		osg_rd_data      : in  std_logic_vector(35 downto 0) := (others => '0'); --              .osg_rd_data
		ram_cs           : out std_logic;                                        --           RAM.cs
		ram_burst_access : out std_logic;                                        --              .burst_access
		ram_burst_size   : out std_logic_vector(3 downto 0);                     --              .burst_size
		ram_address      : out std_logic_vector(23 downto 0);                    --              .address
		ram_wr_en        : out std_logic;                                        --              .wr_en
		ram_wrdata       : out std_logic_vector(31 downto 0);                    --              .wrdata
		ram_rd_en        : out std_logic;                                        --              .rd_en
		ram_rddata       : in  std_logic_vector(31 downto 0) := (others => '0'); --              .rddata
		ram_rddata_valid : in  std_logic                     := '0';             --              .rddata_valid
		ram_busy         : in  std_logic                     := '0';             --              .busy
		ram_available    : in  std_logic                     := '0';             --              .available
		ram_empty        : in  std_logic                     := '0';             --              .empty
		ts_data_valid    : in  std_logic                     := '0';             --            TS.data_valid
		ts_data          : in  std_logic_vector(7 downto 0)  := (others => '0'); --              .data
		ts_data_refclk   : out std_logic;                                        --              .data_refclk
		ts_data_busy     : out std_logic;                                        --              .data_busy
		ts_data_clk      : in  std_logic                     := '0';             --        TS_Clk.clk
		reg_address      : in  std_logic_vector(19 downto 0) := (others => '0'); --  avalon_slave.address
		reg_wr_data      : in  std_logic_vector(31 downto 0) := (others => '0'); --              .writedata
		reg_wr_en        : in  std_logic                     := '0';             --              .write
		reg_chip_en      : in  std_logic                     := '0';             --              .chipselect
		reg_rd_data      : out std_logic_vector(31 downto 0);                    --              .readdata
		reg_cmd_ack      : out std_logic;                                        --              .waitrequest_n
		clock            : in  std_logic                     := '0';             -- cms0041_clock.clk
		reg_irq          : out std_logic;                                        --           irq.irq
		reset_n          : in  std_logic                     := '0'              --       reset_n.reset_n
	);
end entity DVBT2_mod;

architecture rtl of DVBT2_mod is
	component cms0041_wrap is
		generic (
			BUILD_DEVICE_FAMILY          : string  := "ALT_GENERIC";
			CLOCK_FREQUENCY_KHZ          : integer := 100000;
			CLOCK_RIF_FREQUENCY_KHZ      : integer := 100000;
			BUILD_REGBANK_INITIALISATION : integer := 0;
			BUILD_MAX_FFT_SIZE           : integer := 32768;
			BUILD_CRITICAL_FILTER        : integer := 1;
			BUILD_INBAND_EQUALISER       : integer := 0;
			BUILD_FFT_WINDOW             : integer := 0;
			BUILD_FEF_SUPPORT            : integer := 0;
			BUILD_L1ACE_PROCESSOR        : integer := 0;
			BUILD_IDV_ADDR_EXTRACTION    : integer := 0;
			BUILD_P2_BIAS_CELLS          : integer := 0;
			BUILD_SFN_SUPPORT            : integer := 0;
			BUILD_SUPPORTED_PLP_NUM      : integer := 1;
			BUILD_T2ADAPT                : integer := 1;
			BUILD_PCR_SUPPORT            : integer := 1;
			BUILD_CALCULATE_TS_RATE      : integer := 1;
			BUILD_PRBS_PACKETS           : integer := 1;
			BUILD_T2MI                   : integer := 0;
			BUILD_RIF                    : integer := 0;
			BUILD_AD9857_SUPPORT         : integer := 0;
			BUILD_AD9957_SUPPORT         : integer := 0;
			BUILD_AD9789_SUPPORT         : integer := 0;
			BUILD_PAPR                   : integer := 0;
			BUILD_PRE_DISTORT            : integer := 0;
			BUILD_BASE_TO_IF             : integer := 0;
			BUILD_IF_ONLY                : integer := 0;
			BUILD_DAC_PROGRAM            : integer := 0;
			DAC_PROG_CLOCK_FREQUENCY_KHZ : integer := 100000;
			BUILD_PLL_PROGRAM            : integer := 0;
			PLL_PROG_CLOCK_FREQUENCY_KHZ : integer := 100000;
			BUILD_OSG_USE_EXTERNAL_RAM   : integer := 1;
			BUILD_SDRAM_WORD_ADDR_WIDTH  : integer := 24;
			BUILD_CITL_CACHE             : integer := 0;
			BUILD_RAM_TEST_SUPPORT       : integer := 0
		);
		port (
			clock            : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			reg_address      : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			reg_wr_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr_en        : in  std_logic                     := 'X';             -- write
			reg_chip_en      : in  std_logic                     := 'X';             -- chipselect
			reg_rd_data      : out std_logic_vector(31 downto 0);                    -- readdata
			reg_cmd_ack      : out std_logic;                                        -- waitrequest_n
			reg_irq          : out std_logic;                                        -- irq
			ts_data_clk      : in  std_logic                     := 'X';             -- clk
			ts_data_valid    : in  std_logic                     := 'X';             -- export
			ts_data          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			ts_data_refclk   : out std_logic;                                        -- export
			ts_data_busy     : out std_logic;                                        -- export
			ram_cs           : out std_logic;                                        -- export
			ram_burst_access : out std_logic;                                        -- export
			ram_burst_size   : out std_logic_vector(3 downto 0);                     -- export
			ram_address      : out std_logic_vector(23 downto 0);                    -- export
			ram_wr_en        : out std_logic;                                        -- export
			ram_wrdata       : out std_logic_vector(31 downto 0);                    -- export
			ram_rd_en        : out std_logic;                                        -- export
			ram_rddata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			ram_rddata_valid : in  std_logic                     := 'X';             -- export
			ram_busy         : in  std_logic                     := 'X';             -- export
			ram_available    : in  std_logic                     := 'X';             -- export
			ram_empty        : in  std_logic                     := 'X';             -- export
			fft_wr_addr      : out std_logic_vector(18 downto 0);                    -- export
			fft_wr_data      : out std_logic_vector(35 downto 0);                    -- export
			fft_wr_ena       : out std_logic;                                        -- export
			fft_rd_addr      : out std_logic_vector(18 downto 0);                    -- export
			fft_rd_data      : in  std_logic_vector(35 downto 0) := (others => 'X'); -- export
			osg_wr_addr      : out std_logic_vector(18 downto 0);                    -- export
			osg_wr_data      : out std_logic_vector(35 downto 0);                    -- export
			osg_wr_ena       : out std_logic;                                        -- export
			osg_rd_addr      : out std_logic_vector(18 downto 0);                    -- export
			osg_rd_data      : in  std_logic_vector(35 downto 0) := (others => 'X'); -- export
			baseband_i       : out std_logic_vector(13 downto 0);                    -- export
			baseband_q       : out std_logic_vector(13 downto 0);                    -- export
			baseband_valid   : out std_logic                                         -- export
		);
	end component cms0041_wrap;

begin

	dvbt2mod_0 : component cms0041_wrap
		generic map (
			BUILD_DEVICE_FAMILY          => "ALT_GENERIC",
			CLOCK_FREQUENCY_KHZ          => 100000,
			CLOCK_RIF_FREQUENCY_KHZ      => 0,
			BUILD_REGBANK_INITIALISATION => 0,
			BUILD_MAX_FFT_SIZE           => 8192,
			BUILD_CRITICAL_FILTER        => 0,
			BUILD_INBAND_EQUALISER       => 0,
			BUILD_FFT_WINDOW             => 0,
			BUILD_FEF_SUPPORT            => 0,
			BUILD_L1ACE_PROCESSOR        => 0,
			BUILD_IDV_ADDR_EXTRACTION    => 0,
			BUILD_P2_BIAS_CELLS          => 0,
			BUILD_SFN_SUPPORT            => 0,
			BUILD_SUPPORTED_PLP_NUM      => 1,
			BUILD_T2ADAPT                => 1,
			BUILD_PCR_SUPPORT            => 1,
			BUILD_CALCULATE_TS_RATE      => 1,
			BUILD_PRBS_PACKETS           => 1,
			BUILD_T2MI                   => 0,
			BUILD_RIF                    => 0,
			BUILD_AD9857_SUPPORT         => 0,
			BUILD_AD9957_SUPPORT         => 0,
			BUILD_AD9789_SUPPORT         => 0,
			BUILD_PAPR                   => 1,
			BUILD_PRE_DISTORT            => 1,
			BUILD_BASE_TO_IF             => 0,
			BUILD_IF_ONLY                => 0,
			BUILD_DAC_PROGRAM            => 0,
			DAC_PROG_CLOCK_FREQUENCY_KHZ => 100000,
			BUILD_PLL_PROGRAM            => 0,
			PLL_PROG_CLOCK_FREQUENCY_KHZ => 0,
			BUILD_OSG_USE_EXTERNAL_RAM   => 1,
			BUILD_SDRAM_WORD_ADDR_WIDTH  => 24,
			BUILD_CITL_CACHE             => 0,
			BUILD_RAM_TEST_SUPPORT       => 1
		)
		port map (
			clock            => clock,            -- cms0041_clock.clk
			reset_n          => reset_n,          --       reset_n.reset_n
			reg_address      => reg_address,      --  avalon_slave.address
			reg_wr_data      => reg_wr_data,      --              .writedata
			reg_wr_en        => reg_wr_en,        --              .write
			reg_chip_en      => reg_chip_en,      --              .chipselect
			reg_rd_data      => reg_rd_data,      --              .readdata
			reg_cmd_ack      => reg_cmd_ack,      --              .waitrequest_n
			reg_irq          => reg_irq,          --           irq.irq
			ts_data_clk      => ts_data_clk,      --        TS_Clk.clk
			ts_data_valid    => ts_data_valid,    --            TS.export
			ts_data          => ts_data,          --              .export
			ts_data_refclk   => ts_data_refclk,   --              .export
			ts_data_busy     => ts_data_busy,     --              .export
			ram_cs           => ram_cs,           --           RAM.export
			ram_burst_access => ram_burst_access, --              .export
			ram_burst_size   => ram_burst_size,   --              .export
			ram_address      => ram_address,      --              .export
			ram_wr_en        => ram_wr_en,        --              .export
			ram_wrdata       => ram_wrdata,       --              .export
			ram_rd_en        => ram_rd_en,        --              .export
			ram_rddata       => ram_rddata,       --              .export
			ram_rddata_valid => ram_rddata_valid, --              .export
			ram_busy         => ram_busy,         --              .export
			ram_available    => ram_available,    --              .export
			ram_empty        => ram_empty,        --              .export
			fft_wr_addr      => fft_wr_addr,      --           QDR.export
			fft_wr_data      => fft_wr_data,      --              .export
			fft_wr_ena       => fft_wr_ena,       --              .export
			fft_rd_addr      => fft_rd_addr,      --              .export
			fft_rd_data      => fft_rd_data,      --              .export
			osg_wr_addr      => osg_wr_addr,      --              .export
			osg_wr_data      => osg_wr_data,      --              .export
			osg_wr_ena       => osg_wr_ena,       --              .export
			osg_rd_addr      => osg_rd_addr,      --              .export
			osg_rd_data      => osg_rd_data,      --              .export
			baseband_i       => baseband_i,       --      Baseband.export
			baseband_q       => baseband_q,       --              .export
			baseband_valid   => baseband_valid    --              .export
		);

end architecture rtl; -- of DVBT2_mod
