��/  �-�߰B�P��ي�m���+8�KS�����B������+�rz���C�
c�_����b-�����<"��.�� �e��}��oQ۴�8g�%,U�|*-t��������[wL׈]����[��@���(=��x{zRs�f�Cg�н��H���\�_��������U@G[l�Gݹ��W{���ȑ�����	e����Б�䷒5k,���*�'oP�'Fz�q�3�z���XۉERl�"�t�Eޠ��f+�yD�]�X0/���7��l��'��YŌ�=��1���^�9|�r�w�8�#gXN	��@����A�,��A�𞪐j�`XؾG8�S�F�䏬����tZ1I��Z�㓬�c�y}j� ��c~��K��k�\����n�-��[� ���4�"��B�=~����D��-�R���^Ƣ$����Y++�WL2t4?��>��=����,��.��Tt/]x���!;�\��[�x�e\6��،����ج8:۲ߊ�*.ѷ�E��\:Ϸ���1�x*�e�}��0�0��a�5L<���ݮ
r���\.q�6�����Ӝ������9����+�HEh�aE��l�O��:Xұ�U6n�Df ��y�J��� �ij�\�ΧU�א�)+)磳vzV��	�&�Lď�$�n�9@�:t:���O)g,K�[u��yΟ���0�A��;cV�IPK���U�T�L�8m���_�Ą#���U��Β,����3��}��>� ;m�ML\.r��?\��-�z\W[,Q�O�'��=�i�s24�g̈́hP���ʭ��n���Ó�d�ߐf�$������F�=!�\�g�z+&8�|�� �\���C�G@��ج?6�/0�����Dٕ���LTx:(8B��,[9i�����,�;Y d��[5:��d�����y�ݝ�>lmwn~F�%ՈQ8�R�Y�UW�w%<if��R&]��ig ��+F�K�};:� YΈ�\$�U��iEe��޶S���ďk�R'60請����Q�c�@	CV��a�`�����
e�sLdY��)�e��k�G�O;f���/�6.�<�nfCϡ�:2�am�>��f�P���g�Oz��֢����´ܾ��7�1�-��2_ �!8���c�v/��]YK���Z���Y��F�4#�$��)K	�X��Ɗ5�<��]A���0��.r4m��yu�KSOP�N��ݚ-eH"�Z�&!ފ�Y�J���	c��ܾ~�}z�����fS�1�~%���$��+ލZ*�,@�d`�jw'��I�)�u�^�kd�C?#�(b����Ĳ<���p�e�ۍ(\�[P���U Z׼S�]��Ɂ�b�wS�y�]=',B�b��8n^Y�� ��^��O-�%a���[�I����>�`L#,�>��-K���ч���'�aJ�R��c�Wc��3�hX�*��;���~�o�����Kt*��FL�of�_��H�ƣ��}:{T�&S`�ʟƇ�f�M�&��=��B��;c��Z˧�G��=y�a�� ��F�k,�ʝ&�j�5��/+`P�zЗ�s���"��O�?�O�m���;�A˲�*^&9�a	�2ov	cЅ�P���6�ر���u�A�Љ5�����J>�rX�%��YF��"� �Q	������Z�҆v������k�ե�-�ƿ���I���7�V�e�,`�Q�p�|�Y��U��N��C�>�*x�a���Vu�Q�>�P;���]ľ���[� ��N�킈��`����J���AEl��c���^��{Y&{���t ��i�28�-��O[�¹T̹2�PΉ��&����H���p����#,�.&�P��9=`�	=�}88�v�O���P�S�q8�S�6߯5�3�sP�u��O��8���O�5�S{C��J�����Frf?g��$�/*^P�L�'�Z6E}����θ�)���_d�A0
@�+@��kg���.��I7�F����+�Í��i���J�I���?T���>��W�\t��K-�X��m��-�R�H:(�`���8~C�H�3��Y�K���I�|�T����*l_Lz��4R���;�m$����7	_�����G��CR�e>��:�%���T(�U���.�k���W���M%@4���&��Rr���5`["�淃�����'l�;����Ś��#_�Yy�����s�NNR�or9S��T��m��U��fq��9^�5�%��x�1��_�BL�=U�et$�{����=����'��\�̉��#�<�H
�$��0?HS��܊�!��Y�!j.�Nl]S�\�,z���@2����;Y��#�`������+^ �ʁz=	�VʎW�7�5���QK >z*Ӑ^�:�e�`-8�z�$�����;T�A��?��[֨Z6G$�LL�17T	YCj��(Y�D��k�0��M�Q,AN����{s|/��K��(p}�ni��b��H9zkT�T�D���?�\�3��ʲ//�B�aBU�R�]W���'k��moS�n���9�R��#��!��:�ց1�<�J�������E��
�<%S�����-��t�вJ�i0V1�OϱD,g=�����G{�;��!��V1m�������Έ�kK�N�K1O�g��]_c>�6�9ά������@���ң�W����OQ�1vś}�"/K>k!��9�0������T�ϲtvH������ ZKAt��&� ��_p/��`���%т�xs	~�@|����
��!�w?���|W*!x��t�)"`�޶.��eR"��o�j�C}d�c���§�x9�z��?��j7������| 2.�▂�p��>�`�#D�w��Kƨm[~J1h�
U"�}س=������t~;��K��ė�9jlb�>,�-�r�D���˕�@�DJeF�6xsRJ#��%��1Ҍ�䈝d!��~5��B:��7��H��Ü�`�>"�$���d�N�wA4�֖2�]O��VX�`�{���{�3��B&��$g"=|���y��X�#ȏb������o�h��Y���sn\�:_���M/��u�����N��sB�������Bj=m������wo�|?/[Pa�gNm�(���x����=�H �t����a�x����|�m.�ķߓ Q�����5�� .m�(
�O䙯C�|Ðϙ���r���r� z������p'M���'�	��{��i�qT�D 8�Y�Ѓ�:�\f�hDM4�Jػc�O���-N,�A�l�Q�a���ϽA���H���<1�fOx\�����
��;O<1H�e��˺VMO(��*��7������$o�_��"ڳq$��X��p�����JN踎�^��}�c�2��)�Ҕ���ڰ(�+�"�*�nf/H��5�VJy_���ʟ�jԋ�"�޶S�kh��O.ov_��M}0����w������LV�׈��m�U��1�����y�u��P�t�w��@�iV�Y�K>�����t`�aXw��E�5�w-R��R�YL�Oz\w\�ۍ.ؠ���>Tt\<���@E��y��O�s�Ø�6����3��U���G5��In ��~�t�)Lb��,�C�,�#�E�H�p|=�P��P��M�EC����;�	�����i37��W9�� >�)oR�u��9�b�>�Yh4���
�l�r�r������N`�\j?l����+'��ML���n �M2y+3:�=��0�|���a8t���m�ةv��H�G�܂U�	@��%�V�`���b$�J5"�:��H����	�u���VGl�45-����x��̴I+�o��E<m[;'C`�����R����K�G&�FS��� h���JC��疸,WK�9�v�]�:�*u-:���+Y��xmn�f٣��\+qd%��M��?�y,�S��1��Nf�� ����*~��go2��*���r��,�����M����d�
�����$ۜ]q��I��S������Ŭ��V����$�"�u.�Fɳ[=�82�צ���ň1�ެ�Jjc#o9�����s� Q"�*L��	�{"�_�	!o�N2`O�������
���v�8G>�e��}ϻ�u��6���A˝�k]?j1\r�͹s��j�!���s`�O*�M�>z�E��m#b��x�!��@$�]�j���ID��@~fS�>��=!Zݨ�3cJo�}w$��²�1��<�F�켈�����8�ڼ�=32����[��&ˢ���+�ZҪ�%W���-�x�3͹jt����čg��X�F:h|��ޠ���0*�S���m���ٗ�rp��Я��]U[�}�m�d���Cqf�+y1ɣ���$�8ʫ��|v����U�.�H�����:�,���6�h�
�N�c(���v��Xէ2�[��Y�d�W�B;�W̱�)�P��?Е�	�%�oX�v�l�����a/��/ʽJM˥g��L:=�D 4�<x��Ob�l����3��p{2��6��Go�_�t��\�;�D+l!~<1P�H�� ��?�o2��B`�N�	�L�k#50��8��t��=�L|���7�rIo��Ǌ��RU롟l[Ue)lUN�Ё�.��1��݄ytp�z�?k��;���KP���Wh�	1��Z�����2�xg}�N�|-�1�]��$�2?+��	����Z�+�&�c<'R���~_�l��oSZ5y�?5�U� �70��K	��.<#��U� t#$��	�>T4�P���(P'�Ȯ.���H'^��|~"�ޛ�y*�"����?<�vt�B�4���N҈gW$q4����$;�Y�P^^��~^���͕/6Z���o��B��k��0ɖO�ضb���˄�T�Mj��NbdN��/��9t���&�����J�����*V*`�����M&���
�0OJ��q�i�d�v��9#�	�%����mXک��]1����/�y��Y�����){)�3��L�ʪzlֹF�)��*,`�W�4�hd��-����Ə	�k�˨|g�G%y���U�ĉ��։�t�s�6]�������
��S�A!�����!EؤÓQ�6J �5���a�dR�w�<I�&�����+
�=�GI���ގp4�__I���1ƃ�����N�_��eS��*��V�9:0���o����J0�l��_p9�DP�����a����]$ګy�L�4j��;=V����$/�<c:�(>Bӆ�@�J$t�8X������h:^���gg77b销��ǁ��Mn&"��@�Bk@�@J��$>w�ff=%�3 s@��Oj��
bh+H�Ց��+惧�h�g5�FHy����.�y�1����B���Dٵ2=���A0�4��h�݊�3?���!z�R{tNҀ3��x�������y'�0����+&)y����^֣�m.�ܡo���,b��jWj�YiR-���>�>/�dw���
}�$�/�p�����L �q��-,����2����six���mYP7����v��=���ݫ-N+u��2��j]�]��eeGK���t�� 59�V�{�����:J�d9�~7�
���z唡�n��k���"�:��CIo�S��Tt�F�'��x��G����H���oMO�c��V�r�k�F����懶����p^��:	�:>|GI�o�fB.��m�]4.�c:(�WY��zEp�=�2��>�8��_��IAIf�Ƥ>$I36X�[����B���W��U:�ϧk�̑ �4
�F��Q���=�4�=�mR"Q�j/Ym=E��\؎�5���l�,�%S�S�@O_�}��;1�b+��C�҆�%D#�X��&�<Hka��>iiI�x���
H�d����J�I�7�?c�W���U�C4tvl�$�yV��Z���z��/A�(K�3�@�,A���ʈ~�'��A�饮nN_�:�8�[�/��@��I�T��'��zuVu��=���Lq��c�^5��y �Z��� a��R8i{�^�n�,��7r���.mk����1��X:5˸�$질{*U Jcw���F�i�H6y�6ώh�b�JKx(P���%Mqâ�������Z��SɆ�,�U�M[_���f�l�[��R�Ϧ���]�F��3|���rb�*�#�bz+I����;m�0Y�W�H
�nL�փ�d��ѝ
�^gǹ~���m�R�}V�|P�v��S*-7�a�/Wyd�4��v���0��$씪Q����:񼨊���#��7��=l�r�EW��I�-�L��j��l�#�(|�Z����A�l'��lg�e��x�IuX����k�P$�n�3}/qۛ���%MB��A��gB&ɏ��7;fjp&e`&�CM=W)�!���ʦkʥ���W���o`�0{[raZg��{��*n�R�ǯ�y��F^@J]b�\��@ݠ�����%Q<[!Vx��Z���)�h�{�P)��������a���2`!�Ï�]��O9�˺���x��,�����8�;�$��j̨�����EU)Fn�5�!�gc��
+1����y��Zn�'p����x'x���:�K�5W4��yr.�  �� ���钠�/�T;��B���@F����z�/%�p;��5����]38�QFS�}|�՞_^*�����Ŗ�y�?O�{z"��t�^�}H�� 궓t��;E��n��)-ٚS?�X�{4�}��8�`��.^������J	8��.l+4�����Y�(�OAc���#�~�6��fŲ��RQO{K��Wt�9Um��-t���3C��'��u}L��]٫���"[�T��O9�5͵�}׎*��Z��	_(�=�N�=�SM������\�c�0l�{�=-��R2x�a��G�Qiz�E��;�m�I�˴o�q?J^�����u�y|H��'o &#�~C��Olp%˸Ȳ���Vf���%���)>�ޣ�Nj�����0j������4#^��Z�P���y�!���~z��w�45>KM��x�����1��2�di�v����w�0+�	��",ǲ�� �����*�wR�7��}�[w��!Z�f��Bͺ&$h;�e�
6͹����R4���5�����Q�~c�(���E��ā�E��^9�H��9�\��=Q-��/�����{>��$U�Q��P���0��i�F؁AQz]�uF6������]NY54_�ʵx�4	��%�T:�h���V��'�أK�u.k{ǔ!\��@��Eq�@��u�is�ItTu�}5��;�JE�~�r�	P/�����	�ة/WnC$�+�ni��V�,
T����Sx��"��{���[ ����*�<V��*�!'b/�$�D�Gg��N��zEst��i�>g�M�{w얊k��N�IE;�-�T��bn�NNLݐ���Z7tl�W?���+4�Ǐ��Ъ�߂�ڣ���̭�
ݼ��P.�����o�tB�u	�^���a�WMM���S�Ip����5;���P���.���Bf�a���/�4��BU?�F�d	[Yl#��x
o�H�K[Z�Xþ�A)٨F���+�;u�>����ɻ����>�=u����%�[����!2(�O���7��s���adt6�����;��1.��4�cW�Ƅ�0��� ��Q��؋��7�������_ED�m�����è�a^`��yu�9s�S�N.@�Ӛ������:t:����*����cKuA��|]X�/�j�2Zs�*[^����_��Qb������<���<a�����c~T�a���\?�w3Dύ��欩��R:�<A��j�W�R�D(�?V����_Ӌ����,//��.�"����	�e�G���4/C$&��ji<ۀK꛺���Z�������8��-E��B�Ib�"dݗ�_����X�$�6���b��)��a��>�$A �,IK"�C�bQ�S�íu��&z/!�I(GP1��p�W� =��x����n[&.$)}C��b�,�[cn�j��$����ua�g5�ߪ�ڲ���{X�+(ٸ  0�i*,��� ���y���Z氣§��!�����ie�aa�0��z-�d.r����`�0��M��!�YD�vA&'���o�k��+#�-��]��MZ󃭓;�Q^%�uf�c��\h��ї���DYpwiDD�%}���w���B铙!٥�)k�Oۑ�o���8��r�{�#�n��~�W� �tI޻x��n-P��; ��2��g�P�7���^���p*����k��A�?#�� �5Z��_����Wgf�}��h�z!K}N"�Ԍ"��:����bkg�����h��&̊���p$̵��i2��nh"$AK��\����S�)i�e)'̣x;z�{	|�2�2C�B#*�H�犝x�9��4mW��5�]3�X�M} �}άvɧ_h���
E4Hl�"aJ��) ���;�OH�y �Sh��%��9\(�9� ߟf܊.���I�Κ�:$��C��0sK�.���PC�a�W����(Mw����v���O�[�`�3��=1\&$������,J�]��2��S�Ӏ�N	���%"_�aXMң�@~�js�ج��f#�T�cC���i}.	��>~�%zH�)vd�0F�Us���GP�0�&H��)��}T.֌��\)��w����a�KY6c��wF����� �;9��iR&��E�ŋ&ѽM��J9 ���R*�}� IgH�;z��#���Y
�H��(��[y�9�8��������lI���\�$��iC�(�VO��~D��xJ��vl�� ;�1SB|������~[!�(8��T���%���`�k@S��ӧ�7��v��[����m^����k+�������h�m�5,��`2�HѕDN�o���Ci��ﺠP��(î|ڃ6@�C!@� �(�S�E�Nu���ۧ����n��S�+�U�[p������B&��jbu۾��-��s�O�Z�����!�����;Q����=�Q��)<q�yGձ}'�r�����h�_�M((�&��1.������ƪ���oĩ��V�m�6�gb�4�%Lr�&�0h�����UU0
Z��I�Gя�˂:"�ro�t�ϯr�	� �$�.�	6�[G&��H7�p MB���.
�p1AQ૙��x�zK�>�,ONh�6�)��a\'�W��Ý� �!5����q`� �b�_-�:rЅ��M�b� ��@�K�v���XU��$x���&��j�q=���w�!	7���҃ЗAzJ�ݳ��h��T�=9�{m+�Kߢt8@�� q�J������F�Ce��Ԥ�i�8�^����n�j����=x����WUrC�����9uOB��}��e�N%�\J�|%�GѠ�"���&���hQ�����\�Z@���?>OY�{�%��*J��h�[�a��}��R�!�g�r���a���v�eO5]���m~vQ|� J����%�Y�N�|+�-81���jc�V�ew��*��sּ76�ҏ�����M�@��&�?���we>ƩƆ[�������t��6i���T��8
��`��i�/��g8���hF��ʟ8^N��j6����)܌f��镓Hw�Q��z��iK��g�%oc���\�g���aF�����nH�]���$�Ǭ���OJ�B��0�����j'�4�#UAA]���p��B��QmpJy��h�T�+��	��c
29�iu�K71y�4�45g:��L%6Rg)S���@��R�Jx�j�ቐM|%��C�T��.� J�oQu5B[�*VN�G>�ȦB[�v���!�8��/�~k���������Ǚ�i�	��T9J�1��+��(���q��U�'CO���fg�L�M�}�)8��m,܈@��MO��PTVA��mo�ϥg~~q��_��FzZFI�˺C�0�h�F�F9v50���x��8��9w�Ⳋ�ܰ0���H���>����W�Һ�Bg넪p�Q�U��oa0c��Fl�˴����Jb.��	�����L�9����LO�+���ԡ?���߈>�fRTl̰��$����
r�	�����׃a(}���d0yR�eV�*c0ťK�5��A]�o}�>U{���η�D4c���ǀ>P�Ȗ�J�7WtiC�I2}�n؉M ���+ω,�U��N
�d�h3����-D��DW�$�N��z�{]t�������b%Z%�Wb4X�����j�
4�1z� �� u�T������$y��P����������q�i�P��a��؀5x����{��K�˩3(���5=1����_g(����Cq�+�TA���l�x�
5'ϟnxB��?�$F����z����gȽ۸����C�[�VpS����Ԝs�XEX�i�|���OM�.e!�\��=����qTf@9�Q�l�����O�%ʼ��L�5З����`Ge6[W)�.`.����T͋���s�M@�#gV�^�_����)4i�$�T#�d7���2��*�6�$)C����|$��U�V�����ͭ�Pcjj�'�{T��vcAÞ7�����4k���ɒGz�Ӽ �Y��ѧa�z��WLi��W���-�v1w��CdT��ҽ�B�6q2�����)��U-�tY�mn#�Z�U�wj�/��0��Rv�x�����QDK�2�8nʑ
�ʐ�=�V�A���.fEG���wA�����ν��b�D�2lX��m�tzz�(H���\8�#�tv秜1n�5�w�)��,h��]~�t�6�履��%%;�x30�����\�fLS}���#E�qT2���u��w�&#�xe�RsEz샞�R��p��[T�R�Z���
��}F%s����U(�M��]�h�:l�gakaL��=iN=��ĢF��V��QN/�nW�����A�����.1Z�J34�����!�=㷋���S�޾㔳����)���؝"z[X��0|�	Oq#_�I�?y	@c�~u������+-��'g�_`�����h]q��<�-eԭc���&&�Ѥ�f@�5ŭK�˂��Y��	ȾݣN�d�����}�.��!��O�;�?W�)����p�:���m�8�S��O���c�S�����u��ڄ��zS����s��d�6)c� �����ꋨ�F
/�{1golNe�Ԣ��л��)���L�!�Q]�iъw8.���GG�H<c>��k`jW�pfG?��ly-E �����E��p�8�ʫ�fxq'nW+��ls,����X_���v���� ���ו�&��x�`)�-��L��,.�z��&�tpU;k07��O�U���i���G�\cm��>��?�]ߏ���w�"��p�
�M<��4�":n�O��x�2���B�Į���vY7��^M���>����t�у�V�S��ʑ	}�1d^vR����mRN�)z�~\52��)�`ܓu��K��Z�^�y��6M�N����:��'�_S�rNz��^ᰰ��1��|H+�7�<�}��W��D��pXf����F�ʵ�Iȹ�"e�6=P�-R�v[#���%tb� /�=�x՞J�����;�Y@�u�p��ǈ[������ ��@+M���������ս���mg�lz@��í�����Ӂ.��a5pG�A�>.5q��?4̿l���ovwMo���]��TRm*������T�V�R�����7_��́l�k|���:&ى�� �OɤɔVz�|D1�������ȼ�.�S7Ƽ֒2��Jl��%_�Bbඎ-|D�f����w�������۽XH���G��=x��0��>gd�+�燥��{���Y�>�Ws�	B��M�EH��6%?����t��Ri��QU��x�\�^k��:���<xư=�D��_<�p�Ѵ�W䲹�e�TY��i�s{qs�??�r[�D�6���_#8*Mf�s��j�SEE�����;�˄�	c�~oBZ�:E���o'Z�m���z#Z@�N�w���tX�n?�j�yKgI�`��x����~�Ɏ��p��*^��Uއ=��/tl@����@_�؇;�E�eO��n�q�S�4�����.��I��G��He(ۙ�+�C��g/2�~k��0ʃ�����Õ��P��.W��^���@՛�8{,d��\��8��q\W�\�{;����T9��$���b�6�V�'�ڕk�Y�����'Γ��0/�B�ղ6m���7Kb���c�㐜�)�P��N��HY�]%gN��#���/~�����'(Y�EDIU���r���˔���f�f�����wC�ʇ�9Ж����K�磊�^~h�é~�N�a�M�
�c"�$l����^���oA.&��j�ߔҫ'5�Q�wG�T`�g @~ׂ���-MTE=ޏ��.���FjsA�,TT����*�� ����/4E��?Sv#F@܈D�!�!��\��&\3%���(��m�\FH�AP{J1�	�j���"�Y�f��r�����i��m	t�^Ľ"�V="��a�Ʀ&J��F����WȎb�6�4�]�o%d쉗)i���Y�H�� g��%(�X&�[�d��^�O������cҖ��r�*LǓ�[�t�#!Y�&/���X�1�H�\�􇵟L����N��w�/�F���x�P��ga��D[�&��E����.&c����ިAT�F5M�}�2���Ӟ�g�j��Q�q�W�q<�t�Jo(�y���!�]�y"���8��}3�>���]8پu^�L���ù� Od��<�1��%i�;ǿ���+Q���-I��W
+�]_�8���ܚH��O�����a�p[ ������q���01���҆k|��� B2��T��tl�.%D��OC|��+�����g�֌H-�Fᳯ�ܫs��w9fL�>�Ǫ[��/��V��=�Ov��g��R,�)��6�S�W<�ԡ�
�w����ݣb,S^�/p�E7+ �MS[7�٢�.�Jc�Wʬ��������>c~6/uY�-�}��6��gᄥ�o��ϩH�)�zc�����|m�I,4�V~RUJS#Ӄ������/�.�/#��b|ixx��kQ��3��e��eo�k�VV#��e�l����uG�x;K~0�h�_����M�`���A��X;����
��Q��IS�>�b�f����21%gx�"��{t�vt�y	�h<��6BEw�7�w ��>��������ISd�N��{�żf�h}���B��C�9V��DB��T,�n��V,>u`�c}�}�!�-�=��Dq����-�ɛ�?��
�ڟE�K�S��0��`���7c�<�NT,?��7�/2�I[��\� �^7��0ݪZ�<��q�`|�Z69�f#ƕMJ�sb�IY�I������B�ױ��A�󆵁���Iٚ����������-�w�[�ݳ~����p�5�`@��Y�g�K�13��0Z�i��޼+$V"m"�[:�<��J"tWHL%��$�$�AW���,,�8��*��>��tv�9�[b��^N�0nK D\�3��j{�s����Ǌ��E0�;�.����q� =gJ���m�v{�Z���hSH�)��(�sw�?���g��n��y�*B����?��r��13fR��ړ����¤]�Ȑ�x�H=G�r�9�>ŨF)x�vF�=,�Q&�i,��K+�gU���B712��8w���̏6�ҷ:?���h��g��\��Jd5\AE����c ��
r��Y�Yڸ$��T[��$c�&�4�B�\�	�f�e���>*��\�����FY-~���5����*u�w���PCA/e� WG��#[�7�3��ϴ���E�8[IǸR��&�R鹴^�����`�J��s��ga����(�[����-%����6~��S|��`O�k�Bg��v���9����{JW}=�Ë����XX�]�Yv�*���B�.=��Z`���N/EZ��������(�`u'��U�!D��홷V��x����D�3y}j�";�������_4:��˜E�u��l48��Ƈn��J%"9�(�`�����S���\2߿�8�v
��+���j1�<�����)��z ��ӣ�*���Pq������oQ8ڂ�����S��Av_��-N��=3-�8�wk�y/1�p�
������L����Q�ڻvr8����LO��憻5��B<�{���'�)g>1�.�M�:tv���ةZ��}&%|��q�hIs����%5�ao�6 �A%״!̮���Q�U�'�T-ܠ�͆TWЦ��*yȪޢ�����QA�(���2t6����Z�D� ��.��ا�:L���{fb]�`�رm�Hbp+J}C�z~��[?V��
"�O՗����ؿ�j@L�~#���&[��}?�R,�37�(Y����7Kt�i��,��^���Mj	2��R����n�N�a�e�S+�c.�o�S ��@gB��79�E� Mڇ�����`&}��ݞfg�,���v�Ae'h��
pŜQ��^�e��D�aZɝ����_44>"����4��F��������Z�.��o_�	��=v��?�/)�K�!����7i�?c��6�Cj�tCn&��7v��5�P,�J�3Y�"��b�FCL��LU�!��4Pz������|�邦��r�d��x������iC��l�Z�� 0�U�x�iI2���{������7�8��b�=>�۰�Ǽ\��Hk��/����J)3��p�T�(�l:�����W��$�B�>O�3�z�u�uR	�wv`�B�2�sNQ��\��\�Z���6���-]Ո֣�Buz�G��,x	F�7��hK�}��J6��C��_Jz�,3���Vp_y�~ܨ�?D���s�P���;8W�̣��=f_�[M^P�n�"�j�j���r�oӴ�!�g�W�>��B=!?��o���K�X�� =��l�r{P���+c)���"�:f����9{��Y=H�Ӑ�.��n���OJ�+�)�U��3�͕��G�.�b�1gq2A���J�����뇤��Vr��<�����0����H�������d/X�.�
��ٿaI�A������b�a����@�j@�Ϭ{_|�Tr�lU2@��Kt��U�wtjKp���#�ΰ���0�&i�>E�����@!?�=�Y�B%h;�����,@�z�:��f�f��+Q�Buuؖ�dYo�б���Y-�����٣�����]��"^)��=G+�I㮮�mS	��B��nU�D_W�ZT���w�����$A��@c���!�*�gQ��i
�o��)��г^h�ͧ	 �&�� 6*������$2�%A?�*�'��G�S�&�a���!Hl:%\�_�!��6�lUpx��B''���ޓѫ"]aR-Hc(��O�U�6�Kh�X�s&`84�Đ���z�zO��KZ4Gi��q�r�S��Q>�q=p�{�7,�5l�b��]W���G��Z��N/���
��� ��@�἗/#W������F���c6�z����Ky�n�T������v�o�/�����Pr�IF�Eܜ�#¸��ߞu��k�Y�\��3�m��i�����7��� ��漶j�3�C���0��>�΢�8XH�9v��MH퍈=�)��hֱ����S6��tq=ƙu��=��u|O.Q��5�������'�T��F�I1��l�t��&�[�6K��[�^o1�t ��O9n�0O��\.\��T���c�нg���sJѝPy���Yԇ�^� �0�~�Vl�A��u&�"iP��k�c�P�̫�2S~��
$`�x@��C�*h�.>�û��8��=�y�����UTRA��Bcy���g��ΪMi4=&)qM��_�2Q�<	4�9M�u�Q	�:�*G��7��)0��|�4�\M��C�kn�G��DP��Fmfc�G� P�	����G]$q���:���JR��q��N�`�b$!d�k���r�H
b@eީr�|���)�\���3J?���u7J��U���Kn���j
s�fp&±���9K�?;���kK��i�fN�	���o�J�u�J9�[��F����?��i$�I�LkZP����i����;�A�}�Э5�"�)��N��~_� �y��f�y$���c���8�I#��3�Qd�&(�4p��po�A�3�/b���<H�Ǩ=ե��۽�O��s�.B3^I���K��֘ķ4�
MFG��3=W�UF��&w��-q�+񰊣.>ݵ�ӼRv&��̃�Oc`��*Y���æhӊ�<���1�e,bTy?�Ɲ*�`K�iB�8������y	����Q){[b��G���h�M�n�^�8��o���r3�S�Ge�+�H��̗]���>^��N�+�4Q^��3���2�:�?����;${%�x�,AP���](p�����c66�X�0�؇itU��g���
��G}<'����LF��3��n���7��c���2�J��*��T�e�/%S��!�em���y�2�^tl)&}3�rR&�t2Q���!��>�q��u2�#'�4�a-V$<��;-C�S�`p�`V$�]Wu`�4��Dc(����&1ĥ���f����Kg���(<pK�����?��I��_ KX�K������`�I�F9.�#Z�8�D�Ԯ��S�-q�9ٗ��j��������s1X3�f�O�/��� �B[,!\	; >��U�G1.����X���:�ߏe�����>+X��je��h� L�e�2(���*�钔Y�wuD��e/I�R�2��X雘3��[��݌Mq�Θ�̠�Q8��Eqy���tm	�9��;�����#��&��9#��Yl������aŝR�G���P�"�����r�z���'�ft��5H��g?W���G	����B8,�7��˕����0��PzG$Ѡ�ֻ���=�?$�|ДL�Z����+u����.���Ȫ��U�U�C���Q��*�W�q�N�Z��̄�3����-��w�C�ž�"+o-!M�.5\1]̛0�~Ыv�;?���oJ�l��	��v4��_�-O۷�d���0�I_DB�T1�:�(H��k&�d�i��}�zS�
h���F}��}V"�8�q��?LT�-�!7A��<G̬�>�6�n��S�\�N%@���w�F�-/T�
T���]ۦ�B�@�c0S<*;;:�e�^�f�;��!�{J��U�jv��fNf����h��nA��P/�[�;Z�(���?�����t�ޫ��G+����C.�H-�xY������3BS�,��C��;���[>
�k�<[%x[I���Ã1J6+����z�كB[,d�/����i��9�v3��II�_�\T��ݯ��kՇ; E�#� �<Wl�(���9�	�p���{�`0?S�1��nE]��Ѡ�گ�K�;�UL�;�X1�F��r��X���
���t�B}F�L����m۫�f�0�IO�[���2�
���X���]�T�m.��T���Hta�»<�Ѷ1�q�����6�(Fjɮ�>/��L����#DY��;S�l��7�T��1�t�S�\m>�����R��؂j)��c����u�@2!� �<�G�ICDi%�$z�D;�� 6�nBP�r6@=j��-�DfG2-�&�Ճ"kzn�]�xjfs�������'³��M����8�π��H��7���m�@�������.��՞�a�:|�>��w62>��I^r�X�*�$u����)]���D6�"�qq��u��ԇ��+3�s�	Dj����ί.������8��P��[�+4%V�������sJ�����c���
35(��MC�EW����ϊ�V����E�����[�����)�%���݁�A�f7�\��2`���%֊�~ӫx�3�je�:9(p��ǈ�t�?T�(����4ۗ �Q�Wؓ��N���- �|z�1�� �kfk�J
�C�T�U���洐�{�A l�q�i�,z;��������|�V_�ޞ��a-�h�ߖ���q��3PH9��Sf�i7�lm�]R-=��d�2��m!�"��Aa��J���r\��UwO�8��+(4�q!�
��H�����L��#�e���7���?0��P�o�:dL�^�έ`Y$.��zS��U(�f����I;!���iqO����*9��T+�B�܄�������T��W�yvafA}4�O�3��3M�����u��Zf���E()��j �Kዘ��A֢� �9M��Oaw��ӸE�PoB_0��t.�e�_t��/vKK�-ë�I���V�װ�8� �3N�:w��8J���!E��d��&���d�U�@[��&rp�R�o�>�ɉ��d+X�p�>W��M��I��݋՜�ANv<��i�H���d�jHP��܂����ne��)��j���S�iUP�!r<�����fɬ/�G�Ͼ�x|+aw���w��-���3�AH.��S�~1K��x�
Ơ^�O\��P��e;�D���'v��_�w߭�m2���|-���$E] zm����ZE+Ϩ+��L������hEr�Z����~�|�iI�3d���_��m���E%ˑ�]��%�h^�����\�?�0�*�K�x�g�n��k��a�w��7"��1�s�����Q9ZI�����7�/�&�Rv�z��N$�zm����Z����#6�^ VQ�B o ��a������הӒr�q(L��V	����˛G���z~O�ٟR&�����Sq�k��Z���E��+�I��),@zw_��0,�s�,K�N���4 }���xr�,,�F㷝�:/H������B��*ކ�@�f��D��Z�$S�	rTK����,'J� ��Sʙ�0��3����lbY�,�G��� ��x��|�w��v�y��~��*=��	�~�P/�-E��ur1N\�>s��(17�>�R9��v���w���Jz��tu;$s�PG���hS�<��!%���o�ė�J��D�[A�p1�p^1D~:����;���f����َA�!3"h�?79!�P��A��x��~���8c��$},�t=�Am���j�h�P��囧\Q*OJ7���B&ǝ?MID^D8�ׯ����Aq��$k���p�M�+��%n�<�R�^�&m;7=�c�c��4��٥��xB�WUY�у_롎l}F�m��iU;�m��!��@m�$�Hg�\���^-��2���g���u[\�װ���|!Y�Yq�4>��n�!�C@�̴��(LN�ߏ�U��c�����"ԗL�n	�~E2A�@�A'����W�.��c�`�7݄���2!G�+��#�S���ō�k�T9����qWs��D��j�(	��J�I4�>�^��� �Gi/. %ư��S�1�%��puё�������qթ�ftI0aP-��O%���̌68�ؑ����\���`�If�}�CIU3��ldsZ������!���>�PΨ|'���Q$�7Nv)��Kv�#�}=Q�d7��X���!�T�)���R��iyNӔ�Ɛy\K�6=������s�8gޣ�2�5맭�wzF!��3�In6''�q��D�N��;X��j���k�C�����:�r�ww\�xf��:����Vc�`���؝So�h��j�OZ�u,�:08�h$�����r	$OCy9&�_�(�� ���B|NS؝�Բz��.f�k��o�{"�j�Tw=R�2�){��Yҷ�]��`3��J-M��΃�����A�J2O#�-hg�uK�5-��%��"�@�o�|��=0�p��>}K�.�ۚ���gc�ն	@��{N\���b(�|e �ʥZBSc}~J�С��W��I���}G�3W+ ��/՚�D���ܙ<U��} |7�]�x�2��[-W
�-�6K�}0�F��A���ײ�{���>y���<�
���nSş.0]�t�y��R�0s���|�=��}��B����Ƅ;.�J-zV��L��\��|9��Q[��<	�U��0��%�}cM;��zX��MP,�5��:���e�������ç�H��ܪ2?<1/��P�Q:�A���b
5:���a��5��l�}Ωi,�Tgn㠢D�K��!�
����3r�៊�j��`�y2-�Q�&���wh��Q�2�U�c��mG�P�93���f�%K�}�N��!��q���d`ؾV�� 
�N�y�C�怹g��ɮ�.�]Hu�ٜ2���Დ�\��|V@]�2#lLC׽���h~�>R
��_p^L|'�)�6�:(�oC�l�e��-$�v89Sʳ�8a��
w��H@��*�zy5�j�9����{�bL��x�,J#�Gm�Qt"��F�M]s�g�۴u2�	��)1����Ln⥈(:� �.9�o'<�އBw�Gs�f��gY��w���z
ُn�R��T�k�0����+��Z�H6����;�]��wX.��m��;��b���7��S���|j�`�S�y���Esh�
9�O�>��;pTЧ-[�Q��_���	�l=�ޑP�Ꮷ������_ g�!AçP�}�}O���f?��F/�m�َu���q'�سÎ_
L�PB	�_!��+a3�aqq���JI]��8	�ΚN��&��κ��mu@��W;q{h�k��lZJ�kG�����\ﶅ#��X��B>�s�e'�]{T�rH�F%����%�\Y�4dnv�|3I��w��N�� -0�����[15�p�D�o8��n�%��X��. �}IL��<��
�W��u7�ĺpC'�e�R�*1d��W���s�Y:V)��?��R�3��,���4�B���"[��vc9��!ɵ{�R������#�nA&(O��HI)X��qL 侻�
)�z�*TQF��(�|��H����{�S� o@o�]ʅwG�|�VD���Z+��)��XqN/�Q���at�[��,��E)q�Y���Xc��)�R5
}7��OS%(���K1��^�Pu���Cą��N�،��JӇ^��I�� ���rP*gP�@�U�9������-�k�"X�q����3���uM(�fR�\��k+�k��팄M��,i�p�T�_�,�p��Z���ɶ<;��T�eO��F;��_�5 S�p)ևؑ+��p�M���UkH;	z_��D@?u ��`��D���QJ\�V%߶�IXlj<v�W1�d}��(��M��Uo�W��� ��kw֗�e������Z�����٫2mQ�m���,�ۧ;AT���$�ik�;�������� HN��t4��8�d��q�{ۉ%�9�e	c��&\���׬O��}�	R r�{o{��������b@�\�#�P�b�1����i�~풼x�nd�)�v�ǲv�r{`������f2���Fee��4�Hk�)*�B���.X����O���kZǛ�<�/�d�Z{RGzj,�
�^/��h ?�f�����-���ՠ�~%Y��W�u�w9�/~�XĿ!ŻE�-�1���l�c���A����q+e����D�C��p�Mk~�atgxr�3����]���u����Hc=ikk$>�ƶ�dQ�[G�M��ٲ�����!�iZ����>"{�u���آE����F�ƃZ[��d�;�G�W����sv#��&�A/K"�$�)~p"�7�w���E�w����U�Z��p�k�=�՟&���̭�1>D!���0�ƃ�f�1��pL���J�F<��I�d��ߚ�u��2�0�>*H�}�? �Ipm�l�  {�*�smbN�� �\�O�|���K;��&+��s�[+V�a��'�n�|�2ю4[:�����E��+�?s]�2�ݔE�v����FS����m|�KJ�.�f����M?=��.��o�&@ԡ��4����&b� <�)��z�#����U3Ccz���A����,���	���Ҭ/�C$���)��f��:D���k�E��YX`<�� �����
��u����uwMn0:ې_���Z�d�i��}#@O�~N������_q���e�a��@cO�@l1���Y�>�>5y�pY�o�nE�O��޷�z� ���TvB`xAhE �{'�M��mH���#�}�?�
>����r�d�"�(|m�)c6�M�[3*�`������K�*�����T��v�i%��}$ߗ��5��^z�>f0Y�>#�׻�5�`"�D��� ?gnG�o0����hTv��0!�1�>�w�������b�yS�$�� �w�x���<�$a���b6�	u�z=��ma����P�A�(Ŷ#g����JKz}�u.�c�ٶj��B�3_�pD�?TVD�����'FZۤ\�/�d_;�(�� D�ȹi�94h�K�
���Ғ�6e��� wzU�J�� G(kh�n/�Z
ꓩeH")��]����K�Q�W�c��3�4�Q��4	WyO��܈	��-��X�[��>�knm�&�ke����*�_䝤 �9(��0���J�K>�e"4����\o�ka�
�y�U��Wۣ�߹� ���4�	[ꏹne]?��W�$��7A�`@'��v�h������⦛X�@�}7��N�t&��<�1�~�x"�=��Z�K��萯3p���J���d�b\\�7�w��w�þ����:�9\r6tajtU���+\��d�ŋң��n.��z�E�V�g�1�N"�<���o�ph����gZ+�H�C]ćy�k^evv������}�g�4ah�t�JX�d�T�d~�T�� f�Q��C��m��FA|`g��/اϘ0�>*�̯nС	T���^����j����=C@<�&�w��Q�,^��_o��p� ���*���؆њ���U�4� �*S\��Q#�E��y��i��S�WdYI��1�Nsp���9�<�9�͡��W�_��F���d٫^����&��?|Wr�֛W˻x���� ��c`���L�$	%,�ʣ�.Ֆd ����+�����q#��� *�7�e^5�����%~�����eT� �[��kO}�/7?�����GV�[��"�C����A!��)��޹`����>0�QЎ�����=�e�w�i(���p��]��n[�Rs	*0�
���/���#k-jU�� ��A�l�)~�j0�KgF���}�ET)�A��;P}ǻ�"��'���k%O/R�Q���L���p��rӛ���y�Df2�`�AN;ZN�xcW����xF�Ιa���؇��&�3�`��\���1~C�[g�(L� �L��^�oU��UF���Q&�c���Cu9{lz<Ezu0Qq$��v˘m`��~���7"kae�|j�7��b��d��,�q��)>*	į��<exN;��k����W�u1����	=tY@�JٙuW&�{b.�V�-�O����fv���?
����tz��ũ��.VQ�z���>%*�3Ld{�-e����$�-��7?0)?��n�a	�Bw���r��i��g�:#�m�NJ��N�赂�r �#����&�'j���1�[s�����t�%d�6_L� ;YS��� �|V����d���:_�����?��:��)�o�j�Ony�×�Bȅj�u'u�X�������Q ��h��ڲw2ڽ����=)���fBW��q�����6��d�����3#/o>d��K�A#���������Ѡ��@���|s�������A�B�������罏?��E��+�Y4ŗT��ae~��2S9f�-L���X2b5�f���C�.�b�V j��$���l�=a�
Y" �e� ���� ����X�8�p+hl�Ј���7}��� C�( ���1����jw !�K}�#�������hy��Kν���������0�d�!|y��0i[�Y��ୌu)ٟ����Ub���E
J����^�4U�ڃ�$ZL��}�,R��}�b^�	���-͕|� T��>������Hȵ��V���L��4�0��j��<n=s�H�pA.����`I�
����W�}:���g��+v�r� V��V	����y����F����Y��p+����V����쵢����x�K�Ķm�[.�x����{�w+�w��(�A��I)8�fZ� ���U&�%U|~;�
��!,_Sz!�۷�S��y9)Rr\�ǒ��$*yGy�޹�.$��6ӭO;�ߍcl�{e��)��V��+��<�W���R��6����{�
�D��lI�Q�3�.5�� Pk��#��s��V�!  ɋ�����ϒ�a,����X���B�D�Oh�ˉ8�%�=�Md��%��v��mLؤ:2����!t�3yԳ�i	A�܆�!O9��/�~[�ѳT�a�7�����I�ڼ�C��ɂ�B@�a}����
����XoM3q�H���!�/�G�}1��%�Oq�h��ap����T�1�Lv�F���<�<��ƋFe�r�"�kعo�ȋ~79�1�K7����$�Go��
�]5�ܐ3�Xܘ����mT��Yg�(�c����������_Ù�M����j`�X�>���ŀ�4oJ�s���6�7�8��(���6^5��Z(vP���wa��7�R�Ɇ���2y��|�/��=�q��2�!���&�uZ��}�Ҙ�G�5��;A�ꃿ�y�T�%������2�q!�AQB=<��Q�{c��І�S �+4T��\��-H5���DHʶ�rx����kR �b-΢��8H�@���X���[2�}�lXp�3�WB�(����?��&��YQ7B�����e[ky���/�3�i+���#���)'I��lB_t#t�£��P,�[H����w/�5w������SD>?�֛��c�,
�WgL�98ȉ�<|ՌG�7.���.!S�%<����IF�nM}n�D�TC����VˋE�"�n����j�L<�NNE`���Q��4WV3E>~_?<y�a����a6�qJ�A���A�������q3�M��}[F��ĵ���+k�d��6$%��Q�k�ٔ'��8���]Yi؀���8_�c�˸N̢�uf�6e��f�U �Ƨo�&�mHN��yaVT���1��|�ɶ��$:��+@Z���i�B2�������gO��Nc��0�zMv�\�,B��C�y���NlYg����Br�(b'�ϔ�PZ�1��ׁVτr�/�&`���r�c�UJ�,�ژ��3��o�y�˸љkm���	��c�wDW�#]��w:i������������mI��#��1H)!�l<���k��W�U�n�����gUߵ�Ά|�}K��+�mm�t �3E���L˲�s�V�dV0k����y��� ��{O�����𯿠�Y������0�ʬUT��t�U��K4� ���j2��6o�^��,j�8�#0W�\�m�-l[����V���sP��>�x���ѵP�1���J'��#���n�
2���~;_0��Cd%���zεf�dra�a�^yqy �O�q�*� 	�~QpG�D0X8���ͥ!�)����@,�_6��r[�z�,w�lp�Y�U�0��0��d�����b�P%RaV�Yz�xC�\�͟"B��xC�?|}�~Z�����8/�yCnKl�/�	�]<����+3?w�@,�രD����6�)Ѩ,
�\鯖22�5ě$�~��/,���g�V�T���g0��]�ɮ�r�����]d�U�[��d�I:�}���ť���օ�>I^g2N�Za���y�{@�bv��ɸ~������@�e��#��we#��E�����8 j2���;��$��+���c>:yhQ"��������~�)!���#�����F�����W���t��~�=�����m0lEJ��z���5;���ӗ/�S);M��+�����I��8�Ƅ����,Ky�%��g��R��~�(Ȳ,`��d^ ) �K�Tl�?q�ULVx��flc���$�}�]�Zbl헏H�Z�'�������i��H��8I=�`���{RF��]��4�={r���<�O3p������T�K�'sS���7&�/�u�@z9C��-)��}_�OQ�=m�	ee��x{f�I�>�8Y܁y��NC�>���T\\���@.����$�X�"ḛ�	�l�c�\�����Ϻs"��֤�Ş)Gl��QƠcdX���e�v�a�tO۾�1H7��t3�+�	I���͓ė�Q��Xx��1�{��͇ 	I�%��_�'�.^^�<r"IM�F�j��aީ7tc�R$VoV�� �� m'�/f�MEw}�K��hʮ�]�)s��?�� �z�Q��c��|�jmV��@JU6W��?��c0E��g�Ժ4D�֝<U)L0��z���c�L��M��� ��J��n��H��86�k�s��*�H���)�2�(�m���Ob�
���+�CV�!�q�7��U���\������u>%ԇ�|���c��n�v��n+��N�qy��,2d��g���ܑ���.�,;)�UI v�^?(v�HTCbR������UVAH�'�����]
���:;������2�3j�dz��G���È;%1G$x�mj^�I�J�=�{�$��l�k4�[��0$"�\��6(U� d�TeYg%��%���<I��<��fƮ�;nL���r @Vl��1Q�	o���9	��e<�^��^�۩��ڛ�(�g�MI!-2��k�4]U��+D%��_6��"s�3�������L#s��@b�7�&��`�Ƭ�����΂򡨰��B�$CB
I��42�Ђu��R9���L�or����p�����Ecf�Ќ{4��Y`C�r�0'�w(>�H��
0��@���7u�cc2��*���b~D:�V��"��QR�wҘ�C�ma`��? �d2�B��(B�����9bQ�?f�X\�S[xz˛YPhK!�U7`e�����KS;�G�8�O�t��_��k{�'����H>;�f�"1����wr�%� a���� q���'`��b��y,f'� <��:��M�2k�h���x=�kP˰�C-ԌNt�{�Յn�E�-���:^�m�%�yw����-�LO��ߟba�fGd(���9J�������\9q@x�xnA')�d�J�B�hۀlu�{_[:��}+]����z!�|��\�ؒs�=���~�ҳ�7�ZZ>��B��U���c�����e�I�m�ɔ�x�)f�o��A�n`s����~���،�G�=x�r����þ������nh&�Ư>��Į��^�5P�>k�'��m<���D��B-o�������l��Ho���2�;��J��O��� Jc����	��{قk�AG���?>����� �~$�+�y ��D\/���-�}��Y�i�6.c*,T�g��[h�8K��۩��~�������\t�pټQ��#��C5����e��$���m[�\GFk/h*�o�/V��G�tH�ch3s�o���*CCW87���.]�J�]MqKh�lƝX�98@a�i\.���V#����ń{�z��֝�i�
B�@���m6����0�8l97O��yei����MM�5�jTP�*�l.�o$^�]���;�뛡�����"Veʰ��3,ȫ��9�ŭ`��«_��k�IE"2n,;oWQ�<���X�.���$/s�uf��*��Y;h�R�t�m�[~XF�؍/���y�U��ۊ���%��eI��k�������'�Z��7�W|:�d���y	�旽�T6�-��s8��u[�������,�Rڼ��:CAS!;�Ge�����ܯ.���zii��ԭ/��a Z�N:I�7o'�M^A�|�9;A8�u����tW0T��3�q��ͧY�;���rpUq?�$Z�ޘ�c-��19�\,����B\���s�Y'����= �Cj�N6�L��Aي�KK�_����c��Q������ Xy���g�CW�}a=�d%t�n@N��V�浅I�>�{������D�/U�Z��#�D��%��@�L*9�6쩢���_#�rU�׃�?�;t�\�n?�;�;��j����k
n�b�ʸd @�ѩ&�g�>^���Vig�Qt�B���=����
)��+�D/��^���{�d�aw��	�~��~��(��);�F��M&�p��W�Q��)
n`��k��� ����k
ܭ��6oC��\ۛdujY��%����֥��	�ך������Ĳ '~ȸ�b�^A��\����i�pM`�\z�ޢrx��q��X�[C?+.��]��"�MK�\_��Y�lx��g� p��03���Ěu���P��L�Jn���4�LS��@Kx�(�;~��g������,�k�9)��$
3t�cxƴ�JI-M5����.�L/FC������E*�u�G}Z��~��):�� @���c�IM̅�f=h�j�96��q�=�G=�=��x�6!�X��Z���K	����o�F�o�h[�#�?n�����}��R��HCo�{���n���;��U[���5](b��W�10@��f�Z%w��;�A�
VV,�$8eF�^�$������d��~N�(wr�� �ML��x�����|��t鑾�6B`

�1�=@���Ɋ.0����܈���"|��˃�(θO������U�ߘ�%��*�$���F�����'�e���,���P꾝dÖR*$�L��Pȭ�q��`��X�t@lsd�LBo�bgD ��b��@<�U�`�7Z�{ZDYm��T,��]�u�Fa3�����ð	4vcKϾ�G�;�1 Vp�8K��P~�)�9Y^���l��J�+�f��h�����( ���4A����^��B�!��T|��/�T�xl�('�*��`:���k�ū̨���ځ#�e��,\7���J�4#2��Ɯ��Q��*��^I��Փ.�����g���vP�j�Z����q�?��็�B�Z����	P��Τ����:�#� ���wg �>��s�É��q����f�HB5'k1p�_�a+Η&�K�U)����ҟ�  T9�2��K�T�F�r��^Yn`�PS�G��˯x�S}LWmŦ�����0��b�s�!so'5"h�?6�bN������=,��r�p[�Ա�z:�;	.�<�0�;�b��rϫB:�c�.�X]��~�/��AQ��7%X���{T�ŁF��䧠<%^�(��X�	z�ͭ�f�ܤa�`.�9Y�ń�t��[�٦+� ����_�`�*J���%z�����2N.�c�+���Q����?+�O�U0�5��e¦�����s<1�-i�"N(�0�i��@�e���1�����'s�=>!���z�k�O���x ��m8�fv��_��+6|���\*Vu��%bc��|앋�=p��C� ,ZPA�򎱏�<w�"�j�ٜ0>˼�߶��A'�E�l��v���|�C��]�V��
�>m޶��'�,��+6���(ֻտ��t�@ʄ��p����N���Ќ�nE�WB4��!S���]�)ө��U��X!:�:*�#��f�R����]��xp�С�5�msVv�<��MܵX�TM�.x�i����J�a�M���)��)d	�mI�VjN�]kP�����ǄR��r�;�8���d򼲯�{�"@{�mZN]��X7�pu�"�E�L�k�/
����B�:v(ʀ���k;n�?*�/J��6d� $0��3���7f8�~�k�ܫqz7���U����}{IE���r�4 
����߹x�{ks,������V�<�pJR�	
�DӴJ���izq�q������)�ί�>8��g��]`���W��d;M����`�_^C�p��Slj�i=�!Y�C`��qẗ́��h��G�xv桲������Q��h�?����/��A�b��X�աc��Ǒ��Gk����.�Dߊ���gxd�	�͓#�\Ag@�ܺM�U�C�iH�Y�fo���E��~���E�)@��u��^O-�"�7��>��V�3��$�_u���S��2������4b�h6RM ��;+.�~p��g���`s��p�����p����_!��Y�A�ᇧ9t{< ��89�"�� K�r��>�������z��ţ��пT��j
*>*�>���Ɂ���|;�l���\f�A;���03�S���N�K���e|Q#IPl��@&+��N�b	kd~p Bد����Q�Н��7��6gLVxm)#��y=7����T��qv��a����{�E7 ��Cj�O3͓��Ͷ- ��Y���p�sL�<�����7�����g�"���y;�3�=�=��-(���^z��X��r��nt`?#�S�O��.kd�b����S���٪=3�z�sx�Jɗ�~bܰ�lI��]0m S��j����'�~p�X}���Y?<�~;9�z=��3W�_��?$DB�TH�
*15=��׵�j�.��Ǐ_�SE�0�~�&��W-{#��p2G%N�L�=���r��>��mR�]�L�v�h� ��p���,���7�:�-X�W��f�	vQ@c��LG�n���9����b	��CD���g�cST6�T�߁�
�R�{���p�P��Z����#��0ڎl?�%�&�(�	J�����E�e��ͦ����a�f�����ʀ%u��l�hq6�[��~'��3q*�5"�_�K��h]}�En4�����B�-bxQ�N�]��A�k��饨�-`;t&��+k՛Y�a�֝�[w�G ���Q�-p��m�͞!���b����/V_
������C�\JR�>PP�o��CG]⾕��{ۭȗnީ?��� ��ˇ�R�$���AQ����*#O/���w���9����Rt �"NĘՓ�<C�V&�ឩCn�Ĕ:����$�i�� 7 EK�����~�==�M����-	T�'Z�*͟���P!j����O/�k�EK�ho�Q924\b��f�(3�d��RU�㴽�e,c��(ʱ�H"ݕ��׬w��Æ>Y|��=�3�w6�ld��9��̀���|���Q_x4Sɢ�J��xWbn��L�5�#��g�����7���A��(B.��@ ܷ-��9wZ�@A�!;MfA�x|CkM�f��/�z:8�yiu�6�^q�+�}(��P��%�1Dt�E l��"~]-t��yt�B��a�~��d��*oe0�
ߜ��+����[��j*������k/�w̌o�aќ�i�yk<7�ȿ|p��R�)�7�ldR<>�֜ᅻ��pp�i�7���С�����yO��!��HQ&�-"IM������By�J`z��֚!��F2��6�~��l���A���>)`��o�]F�����)祸sлq���a�yn��,`B�:��$�=e�vXW��ٴ��5U�j}|��>�r������|�/H4�23�3J��u;����ͻ�'q���F�EZ5�}��,�G�8��m^\���
���n_�X.��J;f,�C�5���	|�`�X���|APO�E��E���}~D_�`l���5�����׹��|'y��8�wI��O�w��	�y����Occ�p�s��W�;4$H�E������gp(kB���>��gf�m�� (헏����VQn܃���Uq�����M�##�n�a��-���K��=ۤ�	7�b�}�z^T']Pi`chD��Ƭ��׵��&O�]���W{�j���?r���B�U�ۄ�����u�v�a� J:yZ��=���G8������ې�o��qc��Lbjŭ��<<���n�Ƭ�b]�M(��o���nIn����ۨ�d�,ˍL��h�14>l5�w.�T3b��^tLi�H��M�HF8�h*Ċ[���j��vh8�5VD�^��R�x�OWU�|�Le<6�=��`��
˂�~��uc��{:7c�> T�^> ���T1Pwh1�.���jO}��"�s�C�J���L�"w�-;5q��@�u�ϡ�pᰥ��"mn&ϳ�"S`c�:��AszҌ���#���P�>���-z��"�+r�f��di��s$����t��Bp��lK�������ѷ����:0C���A#�`�	)/J0v���B|
s)^�A�r� -3>Sج�
�fmTf�yM9×��#���&�N>��,���(�#'c�����etˣ���.G�m�~���H�m/~z#����e�( #��R���yVˍ'y%a��������'"��l�3E!c�^#s8*>$� b��]�Ӎ�&%�ȩ\)k�eI��m���Y�`�-�_0OBP���ڞ���=*=)d&~20�Ď��*lK�6�/�a!#j���NdM�(�x
�Z�VE���J.�c�)��*
��>�!﶑��Z�/�6?�:��S��B?ϜY ����5���C���I�B�u|�W�U���ʌi&Gu�v�1D,��б/	�Vቍ��d}}��4o������NÓ����D�T�}��®	t�|�2�v��o�7J�R'X.�>r�a�,_�)u��oR��2�;�Z�H8>�4��o�%� -��{VxH`EA;3<*�Ε��\8Q��#s9�V��+Z�ڰ�����_fZ$V�Hg��"L�:�X�7��;�����u��� ?��
^6|$2$Đ���5��������:�q&�"#��n�愛�A>k,��x��V�9?Sh߉w<l��1����^7��I_wvVQ�Vb��Z�Fk��+%�q�ț��@��������ɖ�n��tN+ٹ6��������RJ<���,�l�<S����}�U$� ��&���8mٲ�y��UQ� ȧ���!�V��E�?�{	G,E��Qz�e0�]�QrO%o�B�,�/<�'�l��sb��V�\<Z?��=e&=�E�M�M�A�V����ٓ�k�F�tY7E�%!m���	OQ�Gղ��zK�t�w��f)��\�%�u30����aB�Q����ٽ��	GN���T�7'Inm�(�Vl�X~�	�zn򴢇�����~�M�
�P�7\��0d�C�h��F4�h�M콌N�\s�r���=�I]!M~��SI���B.��[���SM����bԜ�n��q�9�|�>��-;Y5��ʹdE�I *��M��G���hiz�Jۡ�>�3]��7�f�ր6���p	��׆�� �8�bv3�3k���	"�I_��
�m������N��P|9���\pkRb�D�2��\/��3�}�ps��0�D*����]/���:����'��60��s���A�����+�w&�5:�0,�50��nTS�
H`�q]ش ����OVZ��ղ�s�q\��[Ga��W�N+�cfL��ãT��T����p�x"d,�`���E�e���J����@�lH�2פASy�>]0�n�P�ߔ��j�?C��� ܚ���'z#�W���0y2���5:�W�Q�TH���&e���F�R�:�|`� K�ӑU�En�����5�m_0^�ƭ��'�o5=���$y5�G�@#�E'&��W�26h��m͢H���V��Y*0�.����37⫠E1�{bG
��/Ұ��q9�7�}� jGla\�3��X
3��X��R.[���Xu.;?��W(1�oVYдm��[Oہ^,J���M�q�7�=x�f��N��M�����gQ�-�������\xޱ�:������agp��Ӡ-���4�>J��Ԡ^�)�C���a�E���z>N���k��<L�d��n�[��p�����÷��
�ˍ�"Y�k�-Qؤ���/�Ud')<�x��A8�7y������ҽ�������������鶱�k;���S;����i:+��젷VQ���6x.E�yӢHH�@5"J +:8�5Ԕ��
]04�f�F�*���Am���E��-�ѥ�H�^�<����^.�ny�h�L�I�Ɲ)"�dV�>#]�wծ.����j˛����jw�}�HQ�W8:�՛�]>&243NVM�UĲ�����8�hn����W��]�E(1b�B_q[L!B�m<�iMM�!�b�i>�w^���%��-���K�)����PXC��iR�]�D2�e.�2��]fU��N��&�l��c�ֺ����T��&S(?��8U2� ��20�?̼L� �����M��D�V\�������!����.O�*A޿������s��c��g����e��r��i��Q�&̗y���P©N�廬��]��Ɉy�uk_�طٿ�Q�g��2^��|���o��RMh�o��>6�u�_v�".9p��OC��)�-hU>R�q+C����*�o�lr?|6���"�MM���mOK����I���T:����T�:v4�)RL�m��?�3%߿��LA#З{�U�X4��I@^ط�!�����
9�l��7G��8��`�`�P��!�ٖ+WI��_b�Я�Dk�؏��g!����o�=u��wi�kr8��I���*��b7���)q�쁊5��6�ʡ����ަY?,�)D��{�N�&D��Lʚތt�[� ���Qr`�:o_`\�K���Dr�!�=S�;�V}���޹�����^/���u��A!2�jp���w�|у�鑱�h`�����G�a��m�<1��+ƔM]�R�̸ Z�����?]ڵ[H6ئė)��mZ~��=$V;�����3���|���-n�3�^�@ �3pw��4�Χ��8u8�g�ǒ<����p2L�h�n{'��X��p�M�Xz@�������e4g��]��0���)f̵�O��ughn�
�ev�����&�r�_�݄��E���{Ĺ�V��G6�ŞN�<�"l�Yy�gAz���3����F]9��2X��ı5��]k���(#����3���u�l�
��fѪkGz���	�+Ǯ�XZ[|°D��p���P�b��:eR�+�=�'�>#����p�[.#\cb&����I@-n�U���@��� Ȫ\����wq�����O�fx<�SmL���h�}b�Q��w�]Ep�͈����0O AR�rz����}'&ηk��?����EDЩ�V`��S�{�����ϒ�~�ٷF*���(�x�y,�--�{� M�����ߕ�C��Q3�2�e����)h^�*6���Ar�8�"0��6�RJ�֐���q���1i�	i
o�I�j��o>߫��_=�A�|:ED�ɹ?w^2r_�����?Y�I)���k�o�窪�{ �O�?#��O��
x�f��Ţ⩛o@�)!����򗁽	:\ݐ7�F9	2a���J��ەJL��D�֩��#-+�33�����:v�.���-1�����DЖX"�Z�Fc�e��b�!���L#Ώgh`�w���5,/��-�=>�W�4P�*�~c��h�����1E��,�;�埼hS���J��'�b/���r����r'dg�à�ղZ9��EKoVt�Uf��a3�N:a�x����As��Κ��0�[$���v��ƥ�Y �����3Y��}R��/S�:�\7T����*�f_]	?}��G�Or%!���V�}�JXx�۾#a�e㑪����.��)�@�QwoI|׸(0����,�5Q�D|s�[�de����"�꤆� sQ\`��u��cd�H��z�E�9��R�HC#�|�nћ��e�/�')��d�!�Utmv�-��j&�4�]D�QY�h�;��}�hKŮȄ�����ु�ܚi�#2+ڙ�����=���T�7� ��?�_����-������l-��rZ�(PJ��ඪ��*�}E�g�ʄ?/m��2h0� IB>��m�w�X��t�ort�Q�3�����9�f'�M���1�`�N��P&^�}P���ɕ��pf�%���&K�F?!��8$����&����h���x��4�F���F����y�zG1蔐���ԗ�E���H���a������X�
��n�|h����\z�Ѱ��}N��;l�� kޱG���S I�E��(��&�Z��kRƉ��F��}��ʭ�-45*�4��Էh^m<vC�a��"2�A�=��w�)�Y�!y���J��8��A�7��'ݯ"-s�����K)��,CfUa:��L��*���k�t�3�k&��4���#�s����NQ�#t�˔`L���s�P�ND��  M��29ٖ7'i4�s �ft��BA�V?��> �R�'cQ)�r8�V���ϝWr8|�����ha�y!��x��Y�:~��7�Y�ի )3��R���h���j�}���ʼřm?�U�򭖢V�]�ƽ9����D�#�iM�z��vr��|�PW�xBѿ��D�6ί�n�mM���e]`�ѽU�~"ճ�j�n�?0�02T�{���&h��~��T6=�e��ٳ�sǵL�������Kb���9ĹҐ�W����� S|�t��J�Ge�x��ؽ����|]
V��dy ��Xu��Wo�:�X����أ4{��E�)�gγ/w,}�D����L&�C4�i�]ۺ�*(+�W���R�=aL�^���`<r	�x�����ι��z%TQ�}\������a��S֙�+:�ݽYs�i<�]�[k�fw_�t,<}�$���1O���,A���B[.����&{z�p���Qȸ������N��(��[Y4����Y	��U�74,�t9ȮL}n�<JЊ�������t]tE��<��:��,���!�FG�k���+M8�t1(χ*�̅����G���H�ID�s�Ў�R@�=*
��E@V
�ch�C����j�'6������ �� ~[%��$`�� ؙG�|hy��7Փ-fiG��:���x�a�C6��/�m�L��$!�jj��+����v��M����`h��\&�c�3�'�4V��>�-w�ư�W&�Q�>�:�������h������'��]�Ёzn�N%1�4��x_�v���~��z��"��!�� 4�jR��2j
��>���e�1 �9a�K��d59���[>�i) �G���'M[ ry�9>2�d�l�ڂ��	n�0㉀咢�Z�dTB���(�� @,M��o�R��`yK�~�ىB�p��ې�O�ٵ��B���4@tM��D��xg�`�K��~k�hE�t+��=��*{"�F�n��8q�Z��hXOҩ*�xAB;)��K.��~��b:���o��oa�d��'��{$�Gs��%Y�ug�dU��t4 -���ax9�p^�y�R�-n�9�t��Gv9U�Qc%[�'P���;�[�ꎿo�c/&�kP��ԋ�6+�{���S*���M����"Ƥr�?�C��H�N��0���*+�/c�@��~܉U�b.h&��z]�0$CGQ�I^1�J�ࡃM�P9��iޮ>��]�����C,��z1�|�������^Sw��d��U��k8��}t
 ;��sEh���c(����W�����ܜXFɚ�^�B����OO���r������7����m&�₥IENq�Q����<�TR�,�i����'MQ����}���%)��6B��KA�̴2�d�~�Ǭ�$G�"��Ӈ�6L��jP�a%RS�V��I���O"BlG�C?�@k��@P8axU�09�� �nK�b;��F�;�Sv�`3�5g����n(:U����}̧�0j�8jZ���%1�e.rr��7�9�f��榺��ũs��N��A��md\S%Yl���s��1�w9�H�,���j^2�ނ����1��`�}z�w8���x�\�������F��kY�в�a�%_��+�}.�Y���/J��A�h�R�^���f��EbƏ�o<lq'}�9�����t��]xO����������~7��3��$�8��l����m��|9��a�b{��f��OO�#�Sb����Q�b�p�'ʄB5�_��_-�!�3�*���v����@$PМ���Dp��!�\f��4z���	�Ϸ=�o;.3*��.���~��:�2i&��_4p�e�r�H��	��TuD�/���D>��<��ɕ|��%�;��������U���	R���54~Z��u!���-�f�(]�u���{���f��x
��p�j��Tvv'���G�����\A~u�����J��LG�Bl-<���<�ȯ��;!�"������d=�����ȝ��d�@&C���+n�"_���u�>;*��}z?�'>7p9��LP!�X��M�\�{ ���cM�4n`_c�!��65�;.oq��g���f�*O���n;v��`��߲�n��ވ��[�����!VHM��Hud��� ��(��8Z)H/��D2h,u���8�ґ�44k ���2�p�~�\&U}����e�}��Y�`��[�Y��dT��R ���=ÆJ��^x)��x��P4U�����۩�bM��p��:5���S�`,^��W_��0�B����m�LN����1�i�w����GY�����[�]�sg�#�mڠ����:��愿k��ז)����t�S�f7�������h"���o�݀�B����t�ꯧ��4�6�ag[����x�wh9*�%I�������/�ʑͥ�M�eA��������r���eV6�=�-���/ɸ�:`>�<��C�rW���L�\?Q���v/��c�V�v�;��r���/ -'V5+������܁��ê
��9������1�*z\�t�gg.<(�<K���@��[K�2�2�wc	��j¡�?La��ev:�˛���bT
mJ7��{�G�03- W'�۷��4���ny|s�`�8..�����W7�"�<�q=��pkzD����Lޜ^Vtr���]0K2#�������-�1j )�����׬���%K���lԢ��{�����i<�����������Ӻ-�? j*<��۱X�+��e���b�s��^*������zލы"VS���4�r�m���r�Ƚ�|���*����`Q��"R7�V�m&s��	�&���4iʤ�3r�U���� �߽5�}rU����]�S�&5^	ب��ݦ�|�r[�G�^��ig���䱈���������jhUDe����al���H!�E wdiCϘ���B��s�
4Y	af��T�m$_�K搜ҟ���j�s�L�h}^xw�t���U�k���]N�qڂ/-�c�"�����x��.+�v؋�V`��s��Ba�銷',Ϗ�͌ ��=o4>$�ȅ)ǐʳzah�~��{w�E��HF��z�fLN��hJ��|ԬMV���)�]X�R}ڇ�a�2u���I��E�K4����P i�2}��� �f��]��%D�����g��$d4�r�T<#?=�t+Hq��H��2P��h�hJ�+>Ҧs�Cg��_�GG��VW��)d����'QJ��c�`�LąjbT�نG���tc|@(�a�4`��/2��!z��Ig��K�^�d�� �YF$E]s#huj��׀�� ����N�z� �B�G��?vBO��'�<hd{�'��%;�)�K�Yi^j��М �$����^��-)�k���Ќ��!77K~^�,h�[�����79���,�ג}J"V��'^��!��K��b7w:e�FU�Qdt�g�_���"�+�v�կ���&D5H�O�(���\|I�S�JJ�W����;�����+����aɪ�*8���X~^���5��\��rmz[��]�F7+��F��v��x��B|non�_��G
��7I�z���@�[�O
��x���\��0^]l�����<_~Ҏ:/yГN3��o�~5���`0-�t#��e��#�>���c� $�\&�����)K0���sM>�**x8/��,����q�Y�Ѓ�e���	q6����J�^�"��L����W�� z�H���ksu8)�-U%QW�8M:>/�-��m����@�5������'�f�)
��'D ��$�a]�+�hh��BdX�&mҗ���"4Y��a�����0}l�6�Y���9g��7�)��4��o6�o����^�Ӝ�BT I�伦���~BBE�D�S�!}M��J)!j �)��wƌ}v���n�Jh�?;�5�lO_�_O_A�Νp"��R<�%�&@�{�88�ɣ��'K�
�0�~�K�x�*O�s��^��f��T��4㻙*�#��`��w+:���]�.�|{��Y�����L����U�b8 n�p�zlj2\7g�l�ޑ
@�N�/Ϳp�K�B�L}hM�t��)1���,������,Ў�T@�edOlпE	x�U�i�6{^i��w�j#� ��7��Ӕ7����l�u�~鞦,O�#ƚ�D�|���[ܞ�Ap����Q��T�l��[XF�1��]�V[��j�Dѝ/��/V�C�������	�K�{���OL�nĪ�ꫫ�T�e��0��c�? S]����"��������&&�MiM����x:DO��ֳ|���kr:`�7	����Y��>mg�|ޥ|z��-�X[��n�LK�O:����ǽ$�P��(��w�E�sܒ94	Z�@�oA�~Z�=�;Z�łp��E�/9 K;��D��H<s> �����3�&-�N���e4!�e)�|�,����r��>�D)��hSZ����rR��66��]Ɏ�b�_3�X�hq����H��"���cz�[��djC�06�=��z��2}�����6W�*NlF>G>ooq��~Icdd�*�D����d����m��T^����JXA�:'p�����H�Eg�Q�ဟ��	�H~1ӣ��=\�����M^�_*���f�}L��|n �l !��"'$��%75	5��=ϩ�� *�jf9v7:�[O-��u��ͨkʙ� 4�[�\�:�J�1��¬�zE0�(��tMr�O�d}�F��~�;�I���v��C7��ݜ��8m����\�-\j�ҙa���p{��0|޼�c�d�F1�~�����=m���Oؙg�	�W%�eV@#�ڇ�]�����-γ�jۈX4����a	A�8�'3���`dܝKC'�ho<�P�K4��#�D4��Dkf���
y��,���5��40V����Z.�4�+�h�#,�U.�������B�Y߃s�o��W��� ���]��	y�Fp�ԟ�0B����r�15$kQ/��p��ͮ<#�Ud~٢-]���Y�.����4��Y�c�cɯnC	鎩DA�2t�K��bHP��X�5�@��Ҏ���u��4N�sq_�.5��E��	Ct�B�e��#�E�O�����ӟ�Mw�Ļ�GKx�b}{� ����&�����d���SҾj�98PTQ�f����e��9�P!�Ƕ�z�%Rʤkܓ�2�%��q=m�c�hK"�z�'���R�-;���yWt����s��1O.��������%��4���\QN4�z��8ĨP�5�9e9�9^�J�k����[{�A��I��bϤf�H����0Ɵ�Bn�3������d7�����tT�6��A�X�F���Y2Q�Ib{k��Dlʼ|$V�zXEw�!2Z�����{�\�N����;��jn�Bl87_�1fC�S��b|��bX�P4�+�I���kk��}����w�x��Y��
]�⟬��B��]��!v�)c�F�̴��V[�����.%i_� �#Ȃ�;�4`�݄Ѻ��R;�L��QC�GՇT(p���Y�U�x�����S�7RK� 9����Q���d���QQc�WGbj��H���*��E����i��vz�6Xkށqbz�.�#������|�>(�\L��Ga��|��KñS����q��N�3���XQ���T:r��X	eXq_g�b��� 9E/!�o�&�^��?����"8Z�<KJ�������������^����c�D�\U~na2mu�y�L*�!S�ؿU{��7/ҭO��iPZ��-iX���nW�������VSş]tW����I~��V�!��uJ[ ��t��̉���I&�)�!i��պIH�lK�U�Y%��Q���X���U�09�Y��W��.�́Ѹ����vܥ�g�ŢI�Y��t�F)T" YQ�Uk�|��7�<G���\-���G
��{DkZ�D�ܖsj�i!�GC��= ۢD�`�i�1�L�B�C4VV���1����߾ ֞7���A�{c{+���ݮ��ƽ��~�f T���l.�RIꖙ`�3�q[���Q�K��=[�����FR��w�M�-��	M�S���$7	��3#BD����&T�dw1ʂƯj3��8>}
��׵Ԓ�p;��Fu�T,�Z����P�9P����ԣ��:ѥ��z.��A�;	�]|R=���@�;r2QGz��= P��62�J�aNu���U6�G�RS�UD�:�È���!�O�b�"���5�&a� |���0R����C�����l_���;9����sC�Y�h<�-
Fm�`��J���
��à�aP���]_�����I�{8?q�* :��@-3+Q����\�Ρ�8l�x$x�F��!$���$����;��R��VϜ��X���/���H��9���i
���K]�0^�L�ʤ�@���p�Hv���n��~n���B�+*�n�R�ZS�r�F�B
7)�$�䑊�A訥(�t�D�#j��Fն��a�:h)���k�#�,�z�� ä��0'_s��Q�X�c9c�;��3RQ�ʄn�((
=3u�:�̑���ҨI�<��t.^ V՗ܡ����X��SO�~���|)���ل*�_��ޠO��k#2R����V�hs�5��B���C���.���|0'-X�`��\��4�8_����;��@�聱 �uH�� �|;�@��~��3��+S�>�`x&������ǋg?le�D�D-�e޻�!�
���*%��.c��
d�}
0]�l��_p�U��-�.5�z�N�麛�P�>6�M���œ��1C[	�nJ�4Zk���ݻ�1����tV-F)�m��F�����* ���J�v9�v��6�ޞ�����4�މ.���7X���p��*�Q�ʘ�^�p�% �铚�����7��x���&��H��g��F�]9�.����kE�N��v�i���'Pl�6x��e�6A�4�L�38!"��������q,��W���e�&98�$�:-�ʣG�|\��{#��t�h}����)�~�g�vCu��wE��4''w�.CY�~v��-�7���v��~<#��I�ve���]���v�@=E�F��<�TR��3�~�Ѯ�����TUp�� 8mv����1���*9� �	}�E�_r����Km��H��~]GR>Y�jHfNY]�����V
�xa�#�W�̀.[kզ]D>P��پ44���Ϲ�Up�+�2�l`03h�1��Z�
�ZRȻ_�䈂�PH	�/�#��Ч�Ms��RO��ē�z���S��5K~o��,�'���;ҰD
2��(Ͷ�<2Y���7%)B�a��yJ���K`>^�t$�&ey�E/W�:��Q�J/=�����kk���)�sw��.V1�^�d�S�ln��J쿭��`c�@(HXV������ty�.��K��o��F�lx��-��#:ћB� ׵.��!��b�4n����+���e ��.+�DPF�2_��^��1~s�u"���9�2!���v^�̄^�༵|J׶�6U���%�$	ĵh>�%��1�CN�Q�j����Nu3�.��S�v��p����[�Z���V+}�χ/��W��gn���}��n�i��-=V�����E.������?�tBNs"�	Sұ��~Վ��p�UyQc"���� y��:v2�K\d.����1@�$�(p:C���F��(h�S�{TD�kL�D��}�Z,����!q��,R��rà0Y�k���8�y+��	�����t�Q��yo�D�d�~˓jL��S���piv�
2��9�̽�y��^�_Gl%#� ��T�����s���Ol��ds�:�7�,�X��|�m���L������]P�i�Y:�. ʋA������L.�6�:8*b��): p�B�V��ppx�O��4e�H���.�;�b����)Z�N�;�������FP��T�8Y����XtH؂���<����ρ��nB�ӈм�rʸ�� 9�ar�Dj�{� l��k��~�����C��U���y�D���v�"�VT�;�s�Z���U�\*�&s�U��R%Z��c���'`@�L�>�͢���W��C(��Ugz�kbj������� R�dK�:xV���U�����ODJ�YJ�-�<5���!c2���O��(< $I�V�2�I}9����7i"R��ښ�vN���0��L=&v��?-U"��BN�J��V)��Q0�	�G�7Hn���$����r�}dՖ��)ܠ�#7�:>��@CT������TH��f5�5�(�� �&_v�$�."�Y}I�&����_�rd,l�J-P8){N��EQ��ۻ�ż)qօ��V���_�c4�l7�bxpӌڈ�Ȼse+�c� y|U%r�Nj��漽�Dk����.����>m~/k���=��c��zB���ItC����W�Jn���'�kF5_�[�����\u��*��Q 9�<�e=zcI�����Ԗ�����s��gd\���^�t�S���j<�cUF��Ԏ-v>>��^��2� �&r^��<�A������
���-��yl���Qr���0HDm٦m�d�a9U�����a��\O1���'�8��MY�<�H���={v��O���Ƀqw Rw/w�9�;8���>S�?ӳȞ��p�CA)�ٞ���4^�-�2g%!s��M�C�NU�q	j�B�.f�,��WՀʝ��Rn*��2X{e�g�vtL6�� $�>V�x�PX�}�����9k� h�M�~��e��.>h�/�^S�ş#��X�¥�k���L��1��Y��h�h���6�2��"��;!�J����l!)S���G�Б�\��{&�dId-+��������h#�}��r�Ҍɇ�Җ���8��G @�\�{^y���c�!r�V1G����級��F\$UI#�^�
�)��ɍ�y��ԛ/�~T �{�.�T��g��|^�v1r�X����%�#��������e���(B�}�T8����~�%���Jo��ǖ�Xx�r2?lż����lO�	R�TחƎg����j뎎 �u���3(��"�r
��G�tE�:�aT5��w�qf� �W�>��Q�ZiiK���w�]k�".���whOD�0ϣ��5e�}r�~搴C�|?S��5B��&�=�r���R��`-aua�b<�z�"�� ��_�>#�9TFO�p�=aK��t2M��ǃ�P�C6�S���
�{~�m��C�V>���=�y.�I,\#Y_Ӳ�^oȍ�kَP
8h���5)K�t����1��d���+4m��{e�!�zcl�����i���X}��#�WF��r���P��H��m��~��h��U�Kr��ɖ���wJ��JB��� q�� 0��
�u�?�	����B��5��l)�v��� Z�O?�˕���ѥd��y�e[��z����X��,t�e7na|I@jFSM���!�{_]�`g�VqB)}��*qJ���j`�c-�М���`�Z�M4͘��\��I�qKy�P~i�����v���޸�%6�p��qÆRs5��s�s�pFg�{�%{&��>��
�쮫}cxԘV��K�<�+.\T,�@��m5�*Kg4�,F��"}��X+��MA���[�����*�)rg+M*M�@��b�u/�0�1�rg�|������8`%7n�mp�+?���F�n�S��5d�8u�$�"�v��?F�$c����=�����&�қv��m�n��g,�,�ꐠ[�U���;*ǂ���C̞�,L �d.Q2�}�p|1L�o�-�-�_�7�Jo��H'�l	Gd��*^���Ζ"Y#�B6ϑ�J��J6^�\�eF�ů�Sy�DJ��EH�� M���'lx��ݻ�$��uf�S�C�2S�7Tֽt�ujz���<5�l����l�ħ|�V4�H�(�+�o���6_R]�p��^��Hh��/ �K�<��6n�攳�,��	�Ja�ϑW	lhi��Z�����VV�V�F	�9��J�>�Wd�Sģ���P�@'�J��8a���S���PL�دѝё�챿�}��ł��m����ޛ8.�	��{@NǶK�ڮ;1v����y(��u	�m�����o�1S��2���R6xKa�&�Ap��4�겓�$b�v��nq��X		�o���Giw�ݛǒfN�e+��q��NС�a�O�]�����7�%$��r�л���l5�t�>��پ�қ:�3�%	/ҽ}�t�|b��4WK6�0HMb4���e�?�w"���$TF[���R~�?.(�(O�"@u�=G쪇���xz�lp2�����1�E|#�K�Y���k=N�ł�����=@�����̺�7�~�2��X�Ib�	?Ld#�e$]��?����;�!Yh�U=�H��{	�����Ւ�|����%�>4�T!ͅ���Ivx |2[8�0��A�b8֦e��ll��\M����U��K{�ρ�]�¥���"�Rٸw����_�S
9_[	b�������m^���u�}�����*9(-���n��[�� I q�D���3��9F�l�� ~I����rG����{�`�Ew�Q�`�[ o5�l�F��������d4=����?�5/ı��P�uBk�������Ղ���A��7$H�L�k�du��F�����ݗ�njQ[��Y�t|f���խ�����b��N���7.�%1�����/��<��2�1���f�w�n	-O�[ )��
Qx���AROX�e�|Y��g���Ɵ���P���߄}�R��ë�!�T��k�(a��x8rG4 ����3�<�hP*E٧?JFO�9�&�����Z:]X�zHL<|��B�'��,ܘ8�}ǣ�Æ��1�Q���7 �Bm��Ħf	�k�@�}�~47'�_K15�I=��L�Ì0��yU%���g���s�1~T�8u�DA����1gIę$)�;%�U�k�h�W���^�.����o�4�O�a]��s�VĐ�i�Y*�	pJ����A������0=8����~T��;����zD�J�d���M�WZ��px4i�Ie8v�Da�G?@>^IY��B"_٦�\�E:�Y,))����K�y�E�A���鯫v��.h�4o�77圏J�<a��5�(|H�I���4�e�]��kDX��ۼ�{��vħ�C)!�_�6�e�T`J-G71K]�q�v���x��ɣ�Hɬ�+4�
����ǟ���D��H���q]%��]���ID\�=�q�7�{Υ�؄W�n6=�=,bGBO�a�"���a&�Y��Hˊ*h4��Ӷ0�
(G:o�g�In��\%ܛ+#��<��C��L�\�7"uZy�'�M|�������z.÷��N�s��> �}����m�w��a_#3�0H�.��")qk&@\|��e����~>��SnUڧҮL�4WjO��#{:B�H�ۋ4}��D�)�@KQ#��C��|%*�@�������mp���2/ۚ�K��Q3^%ˋ@;�rI�w��U�;i37�f߹08���l��t"��\�O�����̹��@�삂�S�����W�#�D�&�FL3y����<�|����4����s���zK��?Ӳ�s�� �� m
��n�)�����H��CB��pҍ�vY����G_��t�޹��ū���H	��J�e���Y�R�
� ��I�I�QI��qe�D��!dl�h��he>�m��N����\��i����.^ �ؠ�}��	 � 9L�e1>��>�P���΅��{�cu��AT���.ƓS��rn��������Ԧ�g�������ߛc/�9����ᘓv�.������
E&�|	XBi����:�\;Q��Mh�-v�r��gU�H��cb���߄��}VjZF��[�Ο���H�?oX�|����Y�_��.-C,JG�h|J�n�Z*XN�x���j���OW ��ի[��5c����:ތ��F|��o}����/ b<��y�76����y�Ю۲�4��4������� �f ���-�z���֤�̒ā��tܚORw��g�	�&�Թџ>&���b1��k��-�b3C��B�3���(E�h�����V`
J�s0o��V%�x$S���q���0�f�+*�{�00􎫀N�Z'7r�� �<�]�x���Ts�i
X�P3r޵��y���ݓ�Y|���y�Qk	�.i��P�f[2i#�^[+N�����B���~cs��aV��[WRԧN��\�������-z�^0�9��S2�}�T�N���W?J��tr��]�thS�x6�d�����f�)�^)7E����6'�GV��'��o �5�5��;ߨc�o�\�ɵBڑN�E'�����9�kf�NȣB]��w�8��i��
�\��1i�~��^P����s3Fx��A���d�1�U�U�R��\�<d7��Y�#�h��XI�f�R�0<�ז�u'��x����[ï�7��O��)t>�f���ܮ����C�y!/��w-1%�1��l�x!˾N[�T8�a�t�M|7y5T}ǯ��6D�wä�H,��@1��e���əxJ��_<h�`C�l��X��k����-���z�����Z1ՋP��.\=����q���
�j�z]�����X�TF����^ ���#��!�������$L:�*\�;[	]m�ǔ�[#o�R{��B8j@!e� !�L�<�%Sֳ��=Fh��]�?]�̠��3�C����!5K���|��o��ۙ�g"���A���b�h��!��I��|���i1]�[zi?nΨn*$�v�sm�J[r�����g�X�#�n�Xo�W��y�~��h}M�V_T$�vf�CE���	�I�V*<δ~vp.��7��e������47L^��
}
�h�/� )�#u�z�"�&j;������ ƣP�̐�b܃���+����StYЩM"���Q{�b�^�LS�xyx�Y��Jbk��$B������FU�~0n����0~�c�sޫ�VOoY��e��Lh���R��ǆ��|��7-�'�||�-}�dO�nlÌ��-��1�&�c�Y�T�A����J��{􀛚L�����s^t�UM�E^��2ڎ -؊b�>W��|(F4�
rfh0?ɃQ�[��~ ry�-E9G��Xrg��@%�Z�6f<����qR/��)B�>���}��Ϯʢy�g�,���c�����[x����W���D�{��ŮVOu�+x[t�Y`}jLP݀��P{v����V	b�Y�*�I��-�f#��5G�V�C��Z̷!!,�B*��}���Έ���U�
<AA]dȠ��Ъ�IB��vz�/1�;� ���w�%��/�M��0��j�}�I�d,aH��:��	�$������ZYB�p�_{v׿]��	�I+�h] ۻAnߥ4�d3��s�4�>$��Ѳ��L��u󄐘+\�hI�jY)�.�����q5��V������e� 2"Y8oKz�Զ�
�X�@������%����#�ah:Q�G���4��K�W�5�W�!�4/�-�r��B{cs%�*[j�S[�Py�0�xB|�u��������nz�f48�.D#�ߋ�mW���h��gG�K��������$X fȑ�Uv?a�Y�J���"��$g��+U�Cq������J�
"���䭺$���Ձ�J���ˋ�H_P�q ��{bto�0hn�쾒�Jy"�|>#�ѷ�£⥃8�����L-l�/"�h����V�u�g�>����Z��f�P�r���Y� .�NM_~�4���:H�(�/�) �L>���Dr���B��t�Ju�0/nv�E��h��D�(�ߒ����M�G/��֡��\�MZ�%�H�M;�od��r� �W!uK� g�Xg?v��
M�Nƫ��k�2 ��>I��H�sߐ�A1���ᗭ$}���i�5�'4\���;-�$U"VGc�ޡs#��('a�(��s���v>���Re$5d�I�&R�"�0�W�����1A�@�� Ϲ�3ə����'�F`A��FD2'���<�J�o�NdgB�U��+�hj��z�^�/=��Lj�R�D>fG�Y���Z>	T>���R|�x��Ʈl&�W���%����b\>+ _�����Q66������}�� ��M��������j+�v�;�Y����Z��
�����^՛_l�̪_�at�<\I�r#����ΰ���V5�9s�\#f[�~3A�nOH۝[&P�L�-�.���OkwX��B���"x�S.1�:�̾�s�dX��J�"|[�$��ɳ9��!e���Ͳxt���!ک�C)t=��ޥɯ(�c�fuXNa(CML����R�0�ò�Ln��y�a�&=��Ԩ=Z�x�D<���� �ڻ����^��"���MV�^�s[�J�rq�A���I�[G4��d��}�ו���%�NZ3}km����b���ea
�x����t�Kzk��-��0��&˱�]\Pmnࡽmo��I����Z���4�̙v���4mIy&�J�m,�h��[�ny{�)��p��%���2�g�9��Pf�#بmV��h�~T+��?i��2Pݳ�w6IP��~��m�������������1k��1�d���U\��s����$;{y�|�S ���ʞ��)G������� ��&Bk��B���Y��Sr�6�6�`�x��V���'�Թ@qza������6k��Pv�1����!ٚ��GW���ou�V=M���h޾��$�\Ո�4J%�>P�]��akM���ί+�]��j�����@��gx-�#OW�m�!�Vz�j�	�� ��; �_�4t&MC�Z��6�Kv���4;�����뷤���%p��B��GK�0�C����������{�����Tx� .z��X��PSݧ�0�FO�I�JqL���!A�7�	�gT�d��� @���e'd��A���������K-��
6t9#/�B�1Qz�ƴ�]�(���g�U�P;U��V��I��9�R��HX������*�,�����l<"�،H��֫M*��i;Z�=ࠞ�l���Dn1��U��2@[�	=ix�΢;��i���^/�c[�ף��������ʴE3˨I���#2*m����Юpv7�����+l�dɈz�C��\��;o�vp���;^�%�x���M��s�>�<GV��������h��IyL%�V�a�P����A�ɭBm�E��&/���_�řՉ�YSo���
��7ۅ��
�8�G�(��a�0-�4�)��g��)�z�hn�6O=e�bͮ�6{u��(�ّ�9�Y@��n��*�$*KJ�r��H�Ӣ� d�-!��h�����b64dC�
h 5G��l�*���W_lW�a��;�t��ǉ�V7B��A�"��@��Znb���Y1�����z6��:�$��4��՝���e�>����P� |В��X�X$?,�<A��8ڑ��޺t��O��'92�����������G;��FE�nj�d���/�
NUv6�>��3;5����<б&A��1j���qg]��Y�\6�Os�aں�1� �{Q�����ʃ`�eG���PϨ�&�ex�N���s&%�ՍP���nk���F#&��H���4��h�;nU9y�s����Qi9���be6���]�S�{§��:�9`����8$�SӘ�clq4��-)�s�ph����	�џqKTʞC�\�r
R�Q���p��V|�i����(���
ᶜ�~O�!΂�A�
�t��L_��'ƇXx����r�Z�ʍڻ�f� �Z�{X��`���T�� ��cS�bJ����傑�a���k�ޢN|��dW�Z�M1E	<nՓj�*�*��2"�W4�F�S��
C&gK�n����C�D�B�6�y)C�6.~ҫ� z�^})? g�G(��?�);YQH�w���\\�Z{�g[~%<�>��6�=����~��,3@'!��w�I��f�VIÓk��q��e�i3J�J�9c-����-U�̗������3�r���w���\�x�^%�H��q�wR�0q�oO�u��ɸ�m���)��Y��u�S�2�|�Ɏ�֞+%�%����2I9�˂��Pi��Z���|�=p�QQR?UQa<?���z^����Y���ۢp��J
Uʛ(��f�A��m�����I����{fm�L�2�lY�cJ��9�
lx:�`
?H]mA�(�+Z�a��d�W��ES|n��[����ͩn[�8�y��Qj��N��]��N`G��v�[]���GU0/t�H)�d�H�A�6d�8z=�����[���o)���P΅S�7�����Ї�&����F(]���55(�Ws����6�ր6F��[_KV���
'ߙ6�?�
98�_^���X�X���}�p�lV��$���JV�:�����y�j�qN�����2�c0w�*0-
F$!��/e��S���~�#O�,"���I�Ł�{�}��ܧjF�Ls����a����D�Z`���I��"^4����f�|z��B}]�d�8ou\��%!�^��4wO�h�?��!m� ��OR;�6ŊQ��~Ci@�ln��Xv�m;@�4N��L�k�Zod��m}�U
;�Ǚ�`١\����<JL��Wė�#�{r8Jҡ�7��><�׎�Y�4B��5Dώ�F3�����Rm
N� C�O�9S�$���G�<���ݎ��;���C��!1$��uL�g3�)�o���r}˽������'сh}�����i���d��ԁ� �F�E�B������N�e[L���K�����a�,�x2ڦ���e�q��N�������e!%V�%��F�B-����x�O1�2Ah������G<�u�S�q��U�`v@������5�������]GD�E�?s�5�tt�����=� ������eg�$�fH���G�w��Ly��KQ��*����	 �"�"�;�?F/�@�g(�	���:B�u(z�7��+�1�,�%��e!��1��
�����i5:�X��8TH(U�F������:����$[��wn��C��t2c-���5��F͍\���g��]x�R�߲<ɯ��?p�5ۅv�-X��3���?maØ���8�КY楍W����B`���r���T�F��'0N=�����W0��X��W�i���l���]g`I�l�� F���~M��+,�H��Ѩ1=UH<{?�)�ZE��]�REK�cc�ĨlgSz�nV�x�5�a"�ۧ�G� �{��Ӂ=�#�nj��m����a�NF)5���P�W��˨�|p�V��f�>��)s��V�ʎؗ�u߃�o>�A�8QZ�sm䂯6#�̥�][`��d��Mz�"���@�sA�.6�Q � aX���}��^ g|���׭/ܼ��H-�n���J)�fT��{	�V��I�O&n�i���r61K�p.M){��`��E�ز����dt�ߊ"�����\�"5E�����Z}N*��y��u����Ec��]n�7S!g*B*la��N/%�1��YW������,��,�vې��2��\8��S倎Q�{���K�*z@��o���Xtl�P���w5jH��ňpk�1J��Uh9Ϟ_%b/%��k����8Y��%P� 
��.�Q�y�R����_- _l:�Z~U�L��X)A<�����ʠk �Rd�͘��������c�0�j��v1�~�/J�9��-hpH��z���x�DJ��;
��1g���)s�klU5�d�A[�f����y��T}���a�_�R��t�`�&8G���Tz�tg_X�M>:�&zS0$���J�:Q��	�`x��*��e���;'2'��~0�F��C�����އ�� �����,��c�^<�'O�V�Rsi���~nK1�w.A[�c�#g�C�Toºs������٦-{���.����8� 	4؈��R�\��o����B��Ha�9�h��0��"��/��i����A�?���ޭM����-b.���yCѧ���WQ�UI� ě/�O~/��!з,6�>��tgL�(aq����^Q7�&��ÿ�2`�oK<�YG�V}д��&�`�`���;��;՝�N���:����E0M���o6�B�!$B4V��{<O���M�"�{}Y�'?�`��/<�-#��(!t߁�O�9��#D���_�vsu�/U���R'���׏kZ�����[����J��SC�Y�^�vb;%��RI���(F���F�5���o���]u�
60{�i$$�[�f�v
�4lS7����C�Gb~��1f]��rjO��A˨[7�#�Җt������lKa=:��V%������@:�b-G���"U�j��(3��`� J�fPZ�����k�1��F�Z5��1'$	��c�Ŷ"�p���,\��j�ϦX'3�._Y�n~~wr�V�T�$�9�*����cպ���j \�%0��ǉ�ߎ=�BO%�vP=O��]S.���?f�xe"0�JZ��ƭ(�'��Y�;�p�Lf4��Ië��W����x�ҷ4a[��fW��xwa��)7|u0� ��ף�{첶���M��iBh�!����Ñ��{X�Bi'�LZ���H��~��]�o�<E��,y�hEC�BUA;�`o��]���S�DO�ܖ�cQV��N���0o��ک���|�y_L�8@����@@�� ?�M\B7����p֡R�'�V�#^�>�4J<?�F���F�����C���GBSW�9�̿��M0)�cSb�� �\D���D�hJ�<wd4����_��3��9���� �	V�JV�6"��Thx�k{�1*o��(��/(�'	R~�D�=��\�0̡������J��1��р��<�	�c������A��6,<��НX�����]X=E||���WL���f�pػ�RT��圻�X,1�$�D-6���]�m�U��Ҽ��(��
*�=���#��"V��<���~$�|E���?�FT���]��h�$i=�m�KV}D{ ����Cy��u��4qe��'-a��7��lO Ĕǳ�u�.KA&�����M�V��C������b#�c ґY�C|5O�*�d�KVb��Q&��f.�U��ܳȠzL��������Z��ںW����p���1�4ɤJ�.�7�H��,y�0:`mK�l墥�@�����3�@Z˅K�I�N]#w��g(X?�B��Z�N<``/_���r������_�n55�*�v��|��K���׼7/�W�v�Q�5�$/�U�9�Ґ�U|P�r�RֆO���l&"]�ZJ�g~�F�L}��qQ����9���dH�<D��"�4���K� |���	5/�C����rd��
9��Dk+
5��U��7�_s:�lG;�+��3W<M�[[�M,���[�,��>P�jil��;�{��YP������� �X�
�q��Q��u5UA��;�X��h1���:z���~�Z���^Km�{�=�l��(�L������KU'�a�s@T�i�=�~Z�=���,�Ϧ@���n�5��bK�FV�bd=�W~it��D(7��M�'��Vjכ�c�0	o���sN\ ߑ����,f�l%@iD��8۞�Kp�I7Q.��UEAYk(��j�`��L�����ʄ�r��e<��:P:0�BC�{�؂,@x���{���]�� %�
���̷S�g*R�xѹ�-"���gx�	C|�<T��5N���]�a��j.��I��%?�P�0��ؐ� ^aknm޳�҈��+�stƷ�$�rC�-=�a;ʈ�xH�|��u��\�]�-"�d�5џ"�9�<��#�k�Z��a0W��ީ��HW�g�07�bs"-��RP�MZ&�������#�qF97���5� /�gټ�d�ݦ-���Z�K� �J����DRBp�����q�/��_��!�ՠ���r>�et���A��w@���(����N2��	2q丢0d>e�zI�/h�Yo�ez���tG�y?L,����U��D+W*:Xi(&:䋢�NT��u|��I����l[l��F����� -IU��w!ABZK���WgJoi�0L�J���4��s�u���&h~��
|�ն���~��o!26E"�Ն��v{�-�d.P}u���;��9S�@�	�7b�&m�!B���81|z��iB�q���	bb'xFH�d�z'�;ٝ6r�����XvEg��Q�ݿ0ڕ<�g�E͛�����G�y��>>b�P�ة���!uѥ�����ɒ����;o'�1�}�9�ܚ�ya�&>S\���o���0@P��
�@��>��yA�}ƶe���X�NY�����+��k,M�b�[cJ0�Y]B--Z#
Bg_��^�_���q�7*<p�W"w�r��K��0��ҝ�VW�XVH������8��,E��ż��f��2�@������璶k¢��B?�AQ�2�gcs�s�N� �� ��7�^
���Ǔ��Lh���(67���6m��h�J����`��^��D�����"�Gu�A!eD���.pxO��x��P(� �Fw�xy�5^����l���6�k"nm+Y�$i�Yֹ��A��I���1lǍMԇ�;$��������*�! tBGwj���FGm���s6��	�h(Q_�~@�� \�,ϑJ��&:�̂`r����.��.���Rb�r��.�:/�P]	���&��	g5��^3��h�W>��5���b��V5Y7E-�l�Sܴ��6���n���qkaT]PXrYɊ)�]��%L�`�Q���?����s_����mãqŜ6 ��$���D
]<�Q��g6O�>G_����zQ9�;R��숟
ٲ/�R���y;��44��!�WkF�[��}�.���-Y�A�z`1��Z� �
�V
�Eڑ'��y�k)bd�	z&�k���"�qGI�
����{)[*-O���x�� W�sz���q��򪑾��5V�w_,�h�^+r��_�.P������D�5��,��6���Ls�Nh��kS�Ƃ+*@j^�y $R�I�lN��G�O��-����6|[aX}>�8�d���E�F�:�3��@'X�T?ͺf	Ұ=ZY�K���ȋ�n&5��ۿ�R�}V��$. #��<���T՗Xv�zܟP�j���{{��۟��+R�F���N�N���܎K��L�̫��[r�q~���I���R	b�+yLh b��c��U�7�M%�-���fMa'U�إ�K���6�J�����;[}�~R\?���GA��%p�TSZ�i��&=f
��+�t�L�>�&I7�	����Y�m�y��&3�
���L�EL0���S�X�O	�/b�vn_1��v�s:�RK�j4n�kNܼ��a1o'�<о�Q�]�j��U��X�Z�m���x&�~�E1O�=;��oo�Y������L��ʾ�c��1'����=�2��N�H��dLH�	+>�-S\�\�or*�iu�t���$���X�u#���}};\�e�&��ϩ*cM3�R�C	�D�	�`���U�q�*�L@=ͺ�?'fq�_�9>�o=����z�@��K{�T4�o�=a`��Og��
Ȫ^�cEh1�ZX���?Q^뉪�t[m��*���?����vR~_�^������6��Yk�Ki؊������7}���^<�s���+�B}��mjWj����\��?߰Bh�â����gcV|�����k������WGk6��fs�n!H�%�fE7��#�hCz���b��ݝL���kG��R��\V�ڠw�,�gS_�4oM��Ŷ"|�o5[�oֵֿ�o������������ro,h��G���g�W� p�)��A4��� <�QR���$��F��N����TMfVM��B2~�����|C6wx�i��qIHe��%���L'��2G*� ��E#�>�J@�a�C�RU�����oy4(��&��n��^yՓ�Ö�`�$�v�jP5�'ojg���ja�7^?ǎ�� jh���d�nD^Lȯ��:�[qޜ�����y}>m���ڵ�I�C:w��r+��A�ؽ5j��~�=�XB�!�T@H��^ͭ����)�2PD�\2u�d#�ytz��<eɪ�Q���"�1��i�!R>�C\�rDK�������P�,^�3[尽9�[b.�̩6P7<�� ���9!�]o�lzv�D#5�*�F���_�v<�M���W�%Y��s�&��������[�{�TV��"���%˪�'P�ud�	��2���K�!?w\'4p��H�0>h�p�x���iZ��R�z��eΎ,��Y�k�������
KfS�0�P⼰P7%��C��w}k��3:	���7���RG��7Џ���wI�d�U��$�����E�dHPK;7���ʃ)�r\��@�L ��s�4dxTo�:J<���FLv�qlT�B�_p�D��t��YN�w�����i���Y�}[/��	���t��*{*�6���LG���L�p�}�v�*F:�`$�=���k�Wz�7��.�۴>�&@��Y�4 ZK��z��]��n�%8[G�}�#Q�
�JA@�2��	8h*ryS���4���Wz����o~��=.��'PH{z"��6���Jqt����c.�N�lG�,�?NV\b��e�:���$s����ȅE�qH! ŕV�� 7�^�<��gZ�Ҿ����1*'�:�������p�-�6����"EJW641�3�a�E&#��a��٭�������%�<̀s�|O�JmQ�qK�&�#�� �����uMV�.ц[�rc7��$���g/�c�k���R�>�\���m��m�!�.�ʳ�3e���9���\dl�I���h/|tjy��O�����*n�!���0�s<��h2��b"u��0�H��t�x��3��̲uq��v�LW6 ��V���l UYH�8M��m}�����{���'PY.��tˇ��Xo/����D��]�-���JvZ�;����7B��x��P�N��wDp�|S�S/%䖋��;ծ�)ǆϼl|��`�~�{���Lк79p=*fya��/BH����q7���}��j%Ȅ H���$����C�.��;5l��@�R�:;��Jhz�#��M��b���.	�]gi�B�k�z�"�m���7r~�".���S��S<q����4֑�>Q嚹�f��E�B=55�B�o�ơ����J\&B �͊�#_�����&a.Nz���dtA�d��n�����4MMV�`)stde�!���j.=�7E�R�e��{�I��F��'����x�r [�V 6����1�>�6���vn�@"$@Z�+��O����M2��6t	�	~�t;���q��E��y��w������'#�JĠ��j�)(�B�w\R��J����8Vf�V�!��xgۤ�]�*�2�s�,p�$�k Y�^� Eɸ@c�5�V��I��Râ^j��(��.�tn��������T$\�1`�®�������K��:Pk$���דF�t�'
�[�1t1NDa���ň�����N^��b�@����0�g����=�:��	���̻-&q��qA��OY]�Z��օ���nn#��,":{2�z+~|ޢ3�~��S�(g
��6�*��g��uhFm
��Py8��A]Dcy��K���]];�E�J�ђw��Pn'=T�u�p�+N�?��I��Q�'�>wr����s���L�s�f!Bx4��
�@�)�L&���ap��k�{j#gS�p|3O�Ȥ�{��ŅIW�
��q�}��=���!N�ĭz<^o+*"8lE[=Gs4l����-+	5;�;�K߳�-�����;8�)��&�K�Q}$V0y��	 ������ϒ�K,)>C��4g�]�Ad����O�Tyv`q��hy�O�a�~��&z����@锘=o�}����p◄M���|l��U��h�r����V��Oǽ۷�����<�q��f���U*��p~��Xu��<�}Z��K����f�$jGv���%���+��Z�����s*� ��W�F��;��޹� ��HQ�5�U@���2٫��J/,n���_9`�,����wo�~�T����4���j2ցD�IX	^��i/G~�%�_L&�7$N�����♥1�W?����75���n4���*�"�vz�Z9BYw��0	�_d�8j�Ht�QqhZ���d욧5�����;���Xū�	�W�n�mɁXe����w7&���[W�Je��:�/�`�/zK��Kk�V��V�Fdf���ɖ)�rѸ�p�y�T��1^���2��$^����V��q[���+��5o��S�px�.� �03�~Fw,���>��"!��,�Byo�9~^�O�%T��Q)�G�I����{�(/&�;b*W�RD{0�U�l"�`>1%�v���%z����mM���v�Q���g�u`
8�ֳ�aÜ(�[t�xXT�_4�Y�ya����b��N�X�G��C�Pi��W4�̝�����`���f���"%@��h���.�,�TТ�v��o}9��9Ѱ�b��N(����f��٤:�ͳQ1�<�>I�e�}�?�=R�M�:6�JD�4�#��n���G�
Yp���ۃ��s _��B[a��H��x���՘f2t/�����C�Ь�?ڸ���V�Iwڪ�$�f7�b�ƽp)��?���蔤P���%c3���_gA�Ŝ�O:�,C�����[������w��\B}�Pdh�<�g�,g�Nı�W�_5���hϲ��eG�F֋���=��x{�f�(���l���
��̩��BL��G�99��'��P�̴f���P��<�	���t�a���N?AC�i^�D$K����RN�a�恜���
}�b�d�d�8fVD��^��F1�A�t�V��³�Ư�v������֡��,�`\2��lY�O��l�8`��e�֦XΌ���^�G�[���鏳猣/\Ώ�հ1VO(�J��=g\W�b��)��0�!3��)`��(��I������~�mr��>��5P߻��m�V;?�[8�I�����S�n@t�hk���l�Dȩ���q�Lv�L5��6~4]؞�>�g�Z{��~��:�ڤ�{���m�!��*�{�[#|,:%HMҩ�J���!�ai|��b}���05�+Dh�W�f��z
�x�0����sl�J��Z��b��{K�y���C@��%7�!�T���8QX�
,;b/�R�	�<��H������G9q����� ���J��4�~�h�#gpd����!9��6P7z���x0Ы�[��;�*��"k����T���q��x㱲�`"\j��%��YT�rR-����l��y���C�k������=_����L��r`G�87�<�f�|��2�M��)�'dØ<6�	,����++#�R%��z��BȂ�6�l�0�W�f@���_"�1Ę�����E'kN���T>ʬ�"�4ϫ���>���@�xa�U����e��#�"���������	�������l%{���r��5����i�|�z�s������+ը�$�Ŷ�������( �����S,��a�4��P�G�)���$G��.t��Y�Fu5y� �}�)�bd����,��pU����@�V�!�%qWc8B��e���	�Q�Z��3��T�vF#�C�i儖�
y���4m�j	��UWZI��%H�C~m�SkǞ�d���Ыr(����#�k����Lh�oje�4:M�f���K��R��A�0��'^8�^��sC�����	7���N�x� FD��Ҧ0����\����B�ej�O҈[��g��3`�<. 5P�ӌ7<��qOA��s�c��ӧ��#��Q����}�e�Ĥ6p�Yd_tŦ*��evܵ`~���n��M�O�Z-BS�&���P��>cx�L�����A��6�[.�{*���}��9?�ڳ����)r�M���� �xKe��s{�bf݀3wb��ۓ��_hEM�j68O�KN�f����	�d
����PK�m%[jV���	�_{�����UԙV����� �&��&�٬h-��.דJgW�'��kJ��.�N��J�˶�l�q;l�jy��18�	֌8�k�44����U?I�ʺ�=��,Njۥ�W��	�'GoQ���!�\7[|�6�ٖZ�'?H1_��#��#��V�7��!R�F��D!'���63n|���O���o��Y��0���?����5<J���?��e�<�o�Z�u�-UH��y���#��������|@m`��v�wOO숰��mY<1H���㈽\���ȸ��$��R���͏�� Z��+0E�Ţ��D�7R����JG����_����jNRC�ţ��l�:�����a>�@+��FVA���Z��w����5��ӯ��rC��7���En��w[<���N�d�_��ׁ1�,�E��?�Of>�]���v��k�?�����A�)�:��* o(���Y������R�+*���l^R3�l��5�y���I�ń0� ���$�29��������d��NĬ2D��t�7��3�����������>�����3�� 6ij�6�o�KRbIB0��rE/禤 �(��7d��eSɝM5	0��.N�����u��� ���ծ������奲��vk���3$��,^� >n�nm����.Dv�f��u���j�} Z�����#���b'���{9�p�O%����9�8����AѰ�So�%pr�kz��yE0���{���ON�N��g��ƈ�]��J/�O�����͉���U�fv��ϓ���遞����P�z��R�κ��)?U�"OΟ7�V���Q��8˘ҿ2`ҖC+8^=�Z����?��̑n�I�L���5�b T���R��l���Od!P�I����o��$�w\z������K�����x�K�otS@��z�cM��cKp�]��ų�+���k��Bq3%�g#m�iAO�|4U��G�j�ĵ�M;)���T�b�hu��G�w+��CK<_�l���d�Zw���ɫX��ԹKwṐ0z�g�Vd8iNb�b��h*�
θm�$���]����ց��O~R��d�����1�n�}��wF�~��~���%_@Gy�ƽ_!Z0=t6����n"�h:��]>lp�0��VnIi��޾f�=˿[u�#K6h�C2o=��*�%�w/���+���ж'
�F�?����45�J�7kz�T���LY	�&���ʳ�$U G"H������bs	L��P5�R#}EN�kJ��jZ��s�����J�{��l�R�����}jZ��°���!4�YA �=�a":�F�!�z�Y��k�x�gy�Hں%�<ތ����
�IVƩ�?��	z�F�p!�8-jl�n��ꍃ9=��%dꦨR��(i����$>H
�� �Xo��	���T��`��#�BG��@;Iw��EB_49����q����S-�>�Dx&��_�J�s�.'���u�h{�R������aN����X}�a�Kh�~�(�z#c��&}�����w:({���	]�E*5J��;�6��!?�;;���]��GhxH��[�f�5�jȖs���Io.K6�7�v��������$���_p�z�ٔ]�%��!k����{�M��Kl�l�:MF�����3b��X�ަ�V!�)�����*tj�(����AL������W]+�vIt��2c��֕�}=���)�e��'
H�'�l�_�j��C��8�)��D��o�Q�mC�Q]�Cej��]c���ҀV��My����ڋ�|��u#���"pI��5��d���s͍r�ܡl�]��W^u��8�˾�R/����?�>�e�i����J�5���:?�n�1�X�OWdD�&s����\?��$�5v)'��E��;�V�j��{܈�>�Y�'��^G8��p�4�@箎r������_���z{� ٭G:�Z�و��ċ\@q��B������9h��.��	�<��p�`�hs�miv���X��R���:�dKy̳�XV�aRע(�o00,��%�.L7��L��׉�D����Hi�eX�0������#S�ϥg���=�0s�U|l�ҷL+r�;����� P����e�;-+�h��c�(>�$hz �Sa;�yo�K'}zY��#�~l���,�̷�F�պ��Yv���
s�d�~.>C���ۈ~�Ő�7�a}j�3��Z��(4����F߭�����'xq��_�3��B6e��oW��F-7�)��F�F|�L���=�R>�\���w�ՀB2?W��N"PfuyP=�Bx|�)�G�rP���2�MJ{�y�޽��G���M(�~���E��Q�}��N�E؃���6��{M(��ƪw���R�q5����T�"�avi�ì�
�[P*��~��q�o�x�2�1ۖ�;��e ��r_lxz�큑�gEy�6]���34
b�����V�M����7+~� �dK��rY!%�5��� �i%n0S�xsM��q1&�����"�b����-����ˤ�5��ڂ:L�3͛e���ǹ���UB/(���T��"���zE�-ٍ��x�@B����D� OG�����_���.CN�`�6�04L��p���uV��P�,S�нY�K�Wr:�M�L��>:�^W�@ۅ�62�ݘH�vU�߾�� v�V��Vz��-��z{�jr'��zg��J�a�ぷ�= �Q���D�7��QTl%O��i��ذ�����l��Ƈ��Ә��OJ�F��S�LI՝��CplC����}3Bb��]EG�oޅ�*�r!�w�]^F}��������Q��.ن�6l:ջ��5a�!�^RuS��wꞨz#�9M���ɿ�v�$>���j���j�	���+��S�.�2���@��5e�اw��DC��	�B�r��������$3���f.�`�B}�h*V����	8�ۘ8�h*��lh���^��[��ĀX$���wB�7]�=�_I�@���<N���\ԧ���6����n徤D�[7�>ˀ*"W#������������=ۑ�k�������p�^�P��-	�˽��%w���=]X����	��~�%[,�%�'�ez��y!ȏ݅ݰ ;<zX�b��Q�����@<_�5���E�[F|̈���Z�i�`6�'ܺE?1��tW�Ŗ�yGKQ���
8���u��8�
|�`&�霶b�c����,_���Ā�,�x�]�^�.������{$B[Aገ��T=��
����v@�b����gй�j�E���{�G��A`l���)�\��:�K����Uo�f/!�V�ûli�%����'��G�",�W��k�m�=�E���7�,%���z��٦�c%w)�r�L��L	]���0ө`���d�m�����~;�ى�B"wH�~(2zӜy`�q��1��]�Mn윙�d�p����lک�o:Z�̟+�?�H��y4~�S�@/�M��m���v����D�qr@��S	�������?e�xͯ)eo�5j���[�GԞ� �QGWX�!�¾F�4<t�)���X-�L<P!�gE�b�p���bB��{�C_RQ���L6�/���Nb�Xp�V{��������?��<G��C��\�:+�e8�֥���xux|{S�uZ޸�_'gW�pފ��a��+n�j�!�L�3�܋'dǃ�X�Yj�7�
<3s�<����lb��l��'�� z(�h�]�Ƨ =�ylV���cS�3���Pn���S��w�n�ȋ�+�Kh_���G���`��BӉYo��{Z�:��ǚ[J�#dB8���n����Y�H	8��w��1C���ƈw�����y��ѼLo8u�ʓR����oy�m5ESAt��;���x�"��3E�~H�
JB���8�P�q�?Jn�#`nѼ.����(uJ�/�Ҭ�uס�_ꎆ�& C�d�>ӡ3ݥ�#�ע��n���.vƷq]��G�\��/q���D�4�������<����J[��=�߾R�2��\i/��N�?�箊g��]�A����0v�CbL�A�&�h�1�U��� ^.+r��%�<��%����?ݼ�t��!�$��H$�#p���?(Z����?֠4D�`�9oHnS��}'[/T�`@��2�Sa�0R��U.,t�4�Ew,ЮS�9{96��l��ҹ�c�<�@���9.�Y�%�b���D�|-�����Јg�qw���Ќ�զ�7�n��Ԧ!���X,�%�P�%�F��K|�c�<X��xsV<��.u�B�x��̜�h���� Ĥ �6.2�&6-��}-9~�n�t�^��r�|�����g��������+k���W���3������������p�P�i$7�K��!��Y-S���,�P����Q��9��х��?����sZ��HN� �x��z�&.���I�F(���ԩ���؄�)hc�����xݬu��)��l�C_�.2L�bn7᧦�h�o�2�>��
�h��'��p��:/��EH|`̉���d`,c���-Ø��Y�7,R,�j��P�S3+H�=�̶'�,,ʿ��YX��> m=V�A��(�������e�������k��s�G�xM�H�����y�#G̯�\B��Lٌ��~h�� ��D�M�z<�x�EJJ�6�1��{��s@�O0G$*k젒�7{��H�s7���<�#�l�K���UA~�n�@�b �z���C��b�^��^"lMeЌ(eM�g�h#��lp��Z_�����W� �@��!W��6	倩5�'�V�����B/(|Ѧ( ��g���R^X�2�\#9��5h�e��S/�y�1_��G��sr��&Kޗ�1��P����������`K���Y��,��84!v�9�/ ۭc;G�����{5S��r����1%�c�}�9�j� �%�ap{p�5C������������k݁�t��w���:n]���R_}W��_�%\��U�>f>�����Y�gn-Z��:���Hie���L�ú�gu{�+�Z�ǵ�e�>q�f���ԕ6Y>m�D?�㮇G�M�/oI����{K�2��WNo0ޓ{0��c��5J�;�����!fCց��p�y��l�1�I9�^�+7gG��ani�Y���e�8�V���=�]J�U'Z*��w�R�9�xU�j{9��GP��8��3���DcIy�Ɉ+X�{� ���I��ۗ2����ǞA��#4��{�lX�í��莝��GOn+b�P/�^�.�	�]U�eqw�I"�m2����d��V��/OnC��Y.����ʹ�H�w�SW0�r� �z�vc ԠPB2B�e��hP��e폘ӠL��&vkּ3�c�IG���,�3S����o3�ӷI�eW�|�����h*��ܾ��S9IH#�g��DF�[d��E�g,&n�:�.~��i����D����&����������)�<kՉ�<����I�b�6�;��"��\�<hѺ�-v�93�@�k��:� �=&,W�r蠑v�����M͠E؞Sc
�z 8�9H�v�n��I�;��f"|eB�J���c��c��!b_���M��:�Bӧ��A�?�?'M����U�_ƾ����:��Vf���B��3�9�L�������.2g�q��`�����aVy�o*`���:o���GN�w0�𦽫���r�P^���-'�I~��̻*V����%��&�f�gϵ���.�����<^-� �_�j��e��"�%-�>�h��7}?��oA��!,u�@�퍤pw��n��W �!�E���6V��^fS��Z��8Zlrߺ���
P�ᕉ��7(�<�����1�#��Â�G #�8�6g�VmOq�T�ɛ�XN��x��kDk� �M��aT�dN����p1�8�|�X,1�b���d���w��gGc�q�ϳm��7k����(�CS�(_%���ʎ�@�!4O��<����;�3�a�,�;��Z���*�[~��mie���r���^��U����D`t_U{Hs��l�H�
���Ą�k�+֥5�k�=t�/�<�a=��_\Gp�0�dEo����C�d$��eB�.PFL����o~��S�!V��[�*��rڭ �V�A���]9*��\jΜ�q��s�X׮��>.�D�Һ�]�C�32Vsv,�sD�`#�W@����s���Y������jI���lYh���ޗ�o@&IqwǺ����Ok+cT�4��(L��l�
��ԍ!�O�n,�j1��~�s�5�"��ۥ�{���4��D�~X���L���#j�t���ԋn�	�.U�?�g7��V�!���Kuz�O}���=��#�$�����S,^�V�����7��(�9���Q��T*��̱/I�b=�TR�"�ų�a]�~(8;���?d{]I뛟�j#���y���VF�$gA��_KÇ.!�U&- ���\�m�77�y��!&�ΰ�q�L�ҍ7+Tu�	W֍n���m2�	1��<��@��Њ;���gh��� ��FE����}LT��V�0���c�Ƙ����H¡9P���
�~�ʼ�'���WPF�@K��tY�M�Q{
S7l�n��dq�L	H�z��y�0}����P-�#l�(+9��&.ӭ:"a!z���M5��E���+j>@q��NF�a5�8�N3e_-ɀQ��:֌�Ӏ�SAk��ډ�/�[%�n�Zԫ����E&��è\s��`[[�l�d���a;Sf�,�`��������X�W�1>ޙ`��q�2��ȣ��e
ⱥ�{���t���i��m?�% ����J�%̧i֓��g�_���GK������T��_�P�>T�H�6���#��Qr���]vh�2'&���M�P;�C+��8�����ԟ���K|]��C�r٭�
ZɃ�C�̅1�1�h%ji�f>�^/)���t9&��X�l
�Z!����N�X-�u�V��6�>N
�˟i^K���;�0>���{�������<M�ay!h�g(�VpX���Ɂz�eLd��[�=9�����z}羅O��6�C�f�k�9��vn����e�o�N�;���tߏq�6b{��~��&�j ��
�k����qd ح�0ݪ�5pR�u�8����w�6�HA��}r֟�<�V4x��X���/dm 0}b?{�}H�=�%�n�fy������z�_�"�����|\�v39���x�/#��H8�F��>__+x̗	����{Y-
L�����.I��N�3ld�Խ~�VX�V�g���KX�0��ne�p�}��zOۆ������م���֙�h������#�ԧ2�r�F<Ew��4Rv�y�K�i�O�'V�F�2�+�ɡF�O�n#��f�t>�zBUb��ם��k'�D(9x<gL;�L/�g��E+8�{�Jt�ēñ3��L�s�0���hێ`� �^��Y�e�/���B��9nu��x�⨒etCBN���W�Za��q�3�C?�ɗ��Rt}�T� uԌA<!��$����?b���&�+�Љ(\Y_��+����?QKA�I�¿����5�0�r�-OZ�"||}��'���4� ���� �^��9����z�ha�.a(7N�HxQB� <�B�g1)Kqۧ`7Ho������O[D�"��a/�2X��NWr6p�c"[f�p���'�#.j��@��n�w)��]9�Q.N�K������&��__�X9m���t�vF�!�}
qd�nP������H@���/�	�H��1�AR�C��W+:m2?Vn�EXs?�����I�ߟ��4F��D�<�<�Ez�e�B�@�U��R�q��}�mm+b�U���u����!�4�CX1Y=�����7��w���	�`�r��}w�nY��4��<Yq;��<�ގ,=u_��W}��gp*ex�#� l��&⽂ǽЂ�;7',�ydǀ�)�f۟M�v���Af����u���w6�B�z	�V���}��Y{г ��˕�G���=��
{��^�֨E)/y����9���߻j�/W��qg�N����$�e;�%[�!��E&��G�0�Z{�]��6���ycp'\N���`��8C:8�F��w���*I��/k(�T{�����F]�ق����Uхb��4�2�.��8[�Dڐ�+�7[�G����Sn��L�wM\�d~!�S�4+焘��+��Z��EA�n�3�Ȁ��W@-��!T=>F��(�x=�+\��t�$�'S2�#�X8�]@y�Ѭ���Ab�����.��=�"B�d��#GU9ɂ�|����Q]�;�Oz�*�-�T�4�}*r0c�7��I�o�ۤ-�a$�k�I޲��ȧ]Y7bU��6F.�|�4��ƚU�����_����$7����d΍��QU
G	�����.��a&��тʦT�)��� Q�?�
����!�1�H��-u�s`u�|i.f'����H�" EG|��&�x������x���� �,���'}��-7lk����=������Y+5N;Z��Z�#vX�)�&��P�I;����
�i����SƑ5�A仌��h3q`�.
s���-H&���聑��8ȦM��Cf�:Dk'��q�(JY�p\h��l���-TS�)��d�y�aJF�y$��4DZ��ڥ�ù�O�BgI��p�ٛ=�x<E��^-dT_zCJB��w���R������m�"����4g��-�O��%�U9�hbc��a+OǦI���ۀ���tdeמD={An8��Y=�~�
J����*�%T�m���g�4�Syq���|��e<ؖ������C�|��Js�e�#p��U�Sf/d����~�T/�DcOJ����z4 ͡����R6��P&����*��[��0���YӬ�l8ɫ,_N9-�Z�ZZxWC�Р�Wg�$f�u���(S�W&�V�cд]�JB�q�/c�2��;<ӎ��h&�@���.E�j�7r�`({p����! e����+�LdHǊF�&�ĥ��q�'q���e+�x�A%��:���
�_4���g����ͮ�[	wEYܴBIX�#4q�hM��J������>�Z��%@��<i���#%�����>��2���IzIK�+/�qz�����s�S�6t���~��G=&�YM���L�/���ӛ�v,��8��}���b?���{�E	<J	����f��c�W��|�-dֱ�?��%=Q�=4�)�=X�9T�^���*dӛ�9��7w��i��=�F��B&��o���2�� �-���X��o{�($�)_�.#��y���vA��G��Oe%����Q�o�0�"��Û�O|����W6�|��\���kΒ��tʥ����ɞvij(�C�rG)ƶ)��p��`ٙ�z΂��q!�O�z�帴�#�ٗ��0d���%�<߱Ŵn���q� �]�@�H�X�x�j���M�Q��WX����틶�5p?W�Q�)kl&��&�];l��v/m���BD�=%�|�?o8�����/Ǽo�X�2�e0z&xaѤ�+�նkv�d����eI���X�t�A�����JĢ��0���bQI����������>�� �����������*��k��<h��8�S.w��kr�x��vF�z����ƃj�?7;~�3 B�#��-�K�l��a��'~p�X2�֫R���[��!��.��_"�w?���������S����Y���F�|��@`�t4�3���ֻ�i�7N����ˡ5�x��3)L���p���#���D.����8+DK583������W�f�����EW�:�ݻ�p-I����FRcLp�u>�
[�I̮�}�-�m�*Ќ���m!�#�_���1²A���a-B�`�)�k*�R�A'�RU�q����A�Ƹ[9�8����ٵ�T�	U�6<��tɢ�Vǚ80HFpp�Ҹ�n�x� �L���F7k:�VE7����y��M�|c��q,~@�E�3C:�"�V�\a�M�0�rEUj����!b���#n(��S��˝�N&̝�@��RQ��
��:F]�^ų_\� ����Q�s���LqbVV��O�������I����mQ4�ͣa�X:���`�v��!�rCLKy��b@LP�=s�����9q#�O�T�2��H�YՃvcy�	����ɈH���ة�G��l��8��ArRn���ϐ\:��$�G��l��ع-��͔\{k���.g�~P3��8�BFnI�-�����u�����4���\h@�N�;��4�w�z��̟��KM�8����-	)pߎ�_��*;�h����z����Y,�Q�O�({�%��|�!:��:���%5�@��@ ��c��n�q�]y��I��N���a��4w�br�?U�	���U��ewH6j9�ƽO����%���%�n���Jj8.j����EEP���`�`��� PC�Q���UҮ���=��1h2�D�rs}�*�C��Q������JD�{�!�Bw
j/~ZA���8iP��0��G$f9 Q
���2�y�_��t�K�����a�T(}ZE(�al�,xy�a������&0�]Y�'�^m�iӥ�om����W�!7��bf}��a���c��Ss��{�dѢɢ5κ��������֫�R��1�@S�$���c�R��(��l�2<jod ��+���EǲA�^8������xURrP
�Z�$zwFtD�}Ɵ���k�>���\�N_�D^��+����d��n�c��`.�M~6:Jɩ�{(û#�69ե�OY;��:��r3D� zA�7wX�&Ğ�5/z�OW�i�
&���,�pf�`K������X���i ǇF�A2�yB�4u�O�i�.M��f�$1;����5�<�1�6�Gc��~Ը�v�%�K[����~���"X��G
^�������lC�k�=0�xᏽ�d�ojj&_������Y�;cTD��;[󒍍�:W�̡�}�Z��?�44X��t'-8�cb�XX�]ʦ6M�A����h�XW����y���Z)٫��l��$�q��g��a;�ԗ
�x����TH�t�������l�����0R��
9��/�CC}<��� �"q�Ҿ
9�����]�|'����bGK$C�e�A��'H��Q���֗`��E��@!��3&��7ٍ��c�V�>�r2����L��1�^�_�6�)a�m�_���,w�P��}P0�ȡ���D$�Y?-�OL?�����/��C�W&c�	�:�q���`h)h�ʈ�R��dݏ�{�-닺�w*�E��>�:<��Ś��h�����a��P�ܓ�Kl������Vn,NҭB�I��6�.�^t0$j'�ŀ5����^+��
��YD����Y6���{��(��	ٸ7ü�wj"�F�"�ҡ�����A�EW��&O*�7S�@�d߽�X�DO$���q��P'1�>�.m:��?�gk��[�ߕ��B`]P,~9N��h�)��i�
9�����iS�B��ՊN�U�/�+����ueٜ[(]gj�޴��n���Y�#�d]'��!I���Bgۥ��3K� ��4,h��S����̖������!:Ъ���^�⥤ϴ_Yk��J��j̧���"�A���R�K���W\$${����	�4%��d߰y��{j�EEY�䲏$ʍ�N�=+*`.��}�%���9��2g�Q�B_����R�L>̪�j���Q�k��P�]<�GLdT���Z@�(X�-�T��ҦI>M%n>�;�]x1�-O�= <�OjQ���"!�nI��AQ[A)���@��j�a����N�\+b��-��1h3z�dJ=�bA��)p�T��[%
�l��xV�֐��W4�lY0��y���.q*�^]r��'a4[�` ��\}�xY�����!���k��1��ا�[-7
�u�chz�w�`��Đ+��L�k�an�=�e����u
�u�!)C_8�䨅�{d(E�F:�5�hA�|�qJ������]E�3�NH\!�k�D��Z���J"j�i�o=�MGH���?��3�X)8]R����4л��뺩,98�JF��Aj��q�X��"MT��{햷��n��D�"MV�����\�������T4�{Ø�H��ؗK�!=�ba,��iv27�s���E�a5V�ƿ1�J2�~�a�j�E�2�9t�Nɳ�/SK|22�ґ�Q���{�Q��_�(YD��;{`V�{�w5��cߠ�S;oW o22�A|i�o ��z�M�]�������,�&+"�)�e���l6,w�\Q1/qc|�!�b&���A^��	������&�� 	5�4�/t���"����2?���2����vIc��f0�yV�Q\(Z[RMp�pʪ�'�Z�V��$'��b���nN� {��")��a�n3,��z��(Z���+Y~'�mT� ʲ�	�#36u�!C��K������&�4ҕ,�I��!�`�3�nb�� P�ZwP�#�PM��C���D��6�j�r���0�J��6�c���=�=\p�G5"��m�snؤqy+N�����k1Ed����"�Q��	Nv��g2����m���/כ��ԩ��5ld�Y��k!�j �V���Ic��}@+�x��9E�?��ܟ��S��2a+Ee����:�T\4"���ڡUJ��Z�i��9W��(B��[�l��0�N���r�YfG�����%���݊�{�<�Fx=�Q���E�GH8��5�o�~�;.{��[��G���6)Ǐ"���2���He@�h�?�o��\�+����ڲYOiq.,�&�5�	I(�`0�J��0�J�P^yq�%i@09�k���E�p��T�I>&8ž���ˑ�t��i�	o��3�s��Y �åJ|�C�F_F���^Mi~K�ᤥ��Z,q�]Z��"'�k�5?OO��7��6W�W�K���;�"�)(��GHU��(�~�r��J�*���X����YW�����7� X#�u��!�:R��l��l����b�!�����4��YSh��WR����CǙZ��0㻀 &Ah
�%&�]�`�U�Rdox�*��Lp��p��&c`*�����2�	�������ħq�~x&Y�;k�Kx'+gq��uMC�	񞾤J?孏[���}�ry����
Dyrj6w���B����j�OK��E�#�U����
-a��+�|p��Rǎ�C�R�Җ��P}$����3U����ⓗ��^T(����)[RPw�F�@%��P�Z�5�6Ç����B���Q��<}�hښ����qLQ�wQ1��Q#}��s ��,��[�'�x�r-C~�*�ah8�/p���ޙ���N|q�ؓ�W�:�b���A��Jb8U�Й5&T��Fո���KӲY�=�v��.�!|n���CLz�;���c�K,�������봤�J���U�A"]ܮ���M��D#��w`��k�<�n���J�(��]J�㹩D���W�i���EC�D����E�{�-ܔ�cE�����g��Q��"	}{+$�F��|�`�����o����s�Q�{l�r,��53F�_���ʜ�`E��ʫ����%RN��I�ͫ�AO���"'zA'���m9ūR��.�4;۝"�f�\�����rXyPp��9c�=)���e��ʴ���G�Z�G���z~�>�-�>g�+b�=�v!0q�ahq�Z �*�eѝ� Zi;M���^b�o���xwS�݇��8�]1�fSIh*	��JZ������;��u
d�+�亏�OnF&UM0>Y�Zz����p�Ա]m�'�pq3R[S�ZgM.y��~�Ϲ�@�G��~��cɻ����ؚ&�ܷ���6KQ_�uu01�a�+z��zUg6�tiA�	����2�A�~�6�6��n�f!�i*~ɢ̗�䂋�"�Mg�mǳ��W����l���7�t������IM��!��V��E,J?���V�j�z���T*^���c��w��S,(�+���8���R�n��1���Hk���9%�������Lrk�����a:��[������7�c��~��/W$��J,�]�]V�?~n����#)8C@��4�r�^��̚5CN������7��:�T���^k���C�r)��&<N;��T�8��i�RzwsR8 ��KA��EV3�Ò��W�|���!��)��w���F��HU�ϒ,J ��h�A�~T�M~s��C�ж[9��=�U�q�	��74:��T'6�3yׯ`6#�D �4����vnY���=!��ݎ%<��dV���E�[US��`Xs�ݺ�������Ղ:{�����'3�	?=`��sj1�,m�������gJ�WnQ��"r���qg\�kX�`��?_UZj�����Y!�ʃC�QPn��/%
�t���ɋ�W���|�R	��Fl��Jw���a��j)O� CO����0^� Y�i�H�
�b�@3��{�B�D�)�])�Q�5cS�i��	/�0�C��Z��_J����Q����̤�?�$A�DR�u$$iSQ�s�x1���)I�-9uFE�ԉ2�8mn�; N�K��:�8;�Yڕ�J<���!!�4[��%F�k���b=���/��n=��#fr�koQ1�
(R�?�yu���k�oj΀xxf�D�A�Ҁ��jQ��j�<]Ŏ�T�T�X�5��]�pyS�i $�#^��!��=�N��1[G�hY��J�I΋Gv����l)�~�n�J5ܥ�7V錮zz���
++Q���N+���7$�6�z����eĆƗvQ���0�ʧ�#�:�iA�;��	JI��>��ͥ�dbܺn1���5��Ȑ�*�M@As��mJ���?4̲���;�(!xjF&�x>�	=�?R$Ts���`ä��3�n#��ӑC���E&o_0��O�K�>�BU� `�����z��Q5V�]�T��-h��Ӌt[��o��a@sn�_��&G;�;�����HtuDG��f�\������t ��1C��L�D��6ۦ&o�b=+��q!B/����M!>+�)!v�{�g>�߱�H�:k��k���,\�ar-�Js[f�z�������2�>�H�*ݠjIg^@�Yt�8e���%��/0�-�ذ�L}ypG�UK�q�������M���5��\�YD��?�ׄ��s7��ɺ�WdI&�ߩ����쒹2OgY����|�/Bǌ���R�pl���xM2R�H��vuXN��Ձ#�5��e�r��
O���#L�}|�2�gE~��y����"��SU?S��3�6��Ͷ��$9�>^ #����>}"��+r>i���a���b��@_D��?#�&�p�#�MRY*��jE���Ʌi�������L����;W?�?J��-8�T��w*=Y�����_x�3��l�>�̎�u�Λ�▘����Q�B�	,J�mK��E��|�����0mmK:�?��%o�H��rHӊ��U"�	\;��9'���ێj��Z$�:3nW��A,=���J�����*�rۚ�Q/XO6�A�����*�񌚢I�"L
�W����+�lNc8��0
��09���[V���:KRM�Mk��T,��b�.�j��h�B`C-uQ>Ķ�!�� T���,����E���Ц4��K{�'��R	S��W��k��}� J��zm����㿷�K��l�􉮨����!�_{vB�yl�����/A׮��/�iƜ7'�b2���o�Ԧ����4{1�Яh'��l�SK�֕r�.�Tލ��O�̈�1��z QB������b����j_��4��={��Kx�Ĕ}���9�Q�m�Y%�ٙ7�Qi\���I&4*���j|��)�n��ݡ?��x�Y����ߪ�Ҿ#�.O*Z2�W������a���Di��}2����Fa��T�pW���g%���	I�ߘyZ-�����>��$m�s+��#U� |��0���ܰԲQ�"v'#�iB�A���AA Q�ߔ�uA0)�ɹ#��:�Gd����r;�`�������&#}�b�t�X8#�C᭐�n���)/H)���H�E���� :���`�Ӻ�� �*�*C�o*fDT����'Σ(k�p�}+���-F��/�m��T�L����1�r5Y%*dͲ&��K�~�
u}��LQI����n8�WJp�4K^j�ͦoe�}bo�����S����X�vX<���\�3�8�G��aH��@Zn�KWl�����2vJ�5��E�O�?�[�D.UYC�^\���-9W�JS�Q�U����5A���"�[�7���vG-I�"�ƈ2�fQ޾<U��iǛ&zcD]�Ka�燤e��`�B*�����vӫ����>.�t���2�@�RF�DK~).	�h�-P�ӡ���������Tv��9�z����P�wǼU���i�>�v^�O�>�Skd�OK����ܣapVq�e��,cJn�F��=YR�%�n�@(-3ye���}h�~OƄ���%�I� ��S���Υ)B�3��F٠i���ǵ��8ЙD����F�~�'�&��)��*��+� ��E(�O��u�T�������i���M4+�S��6]{�)�y��{��
�<�oǶ�.��v��R�V�Q(@������"g����h+ْ��-G2Yx7���
7 yB�� i�y�u����ed�Q(Ԁ3��r#���<��x�
�|��E�B��0:��ܖzaJ�R�Bu��`v�+v��[�ZdI�2�tH�P��Y�=�V�$��?����/��Q�ьD��z�**T�������*�¾#�R�`�M�'����_�l�-�V|x�� D���^�P�B�+������� �V��{�P-8�Q�n��u`��Kڎ���g�|�5N}�Ĕ0� �K�|��3|'����?��b"0�tu�-dX��P�\��\ ���%��=��7�g�?���+V��5S]�XmI�[��ؕk��#�{�Ƹϸ}P�\���!c���Y��}���1��Z�0�Z���;mP��1Rhd��8]UmB�	T���z����=�h�־zk�!��$T�j�jX�M�zi.R��x�{	��_Eb~JdWT�.?�fM��6�(lf(�l���tu���BV�MT~��k�g?ֈ��;$Y�ȓ`w(�%6�p��9��ы�?#���D	��-�bg<Xn�T{�dpj�� ��VBK�۹�܅(�m82�t�h��6�(.��:�� f��b<��������D�p��ۧ�141�'d��6z��F̢�|�(*���:n��TRN���M$���k��r7z�MQ�.3�����Lzvb{�(�r�@�e�S]¶�Qa*���\����{I����hs֧��J�rb s���h�B!�뫷��Z\߿������
!�O��&����I&ץ+�vĬn�Uz8��T��.k1�j?a��GE�~Ǫ����}KC��-

W�i�v�i�#�A���*�O5����H�#cߢ������C6�,o�V�ܫ��:�����/��w�[�P��%E�q$xG�M�����悙�O��Ku餕F}��	T1�I%��T��?�Y����2��Af8�o4����pD='F��o/��`�9�B�_C��UMg��蚨k�2x��Nm�q�q�/ޮ��[xU��HMU�6��F�����41�t��
T�Jr�R>8��ޓ�K��m��W{�N�Cɳ�^#�(��@�o�1���n �'@�ގy2Vv�'�BA�@��zn*�DԑpbS({vpEZ�l3�_�a�Cq�>�օ��E��Ad.X���� .����67����!���x#�;�TN�)+�X�������:&�%�z��������AQ>���V����	}3��EeHx`b��P�s�/kB�c3/�rb&��>��_�p���Q!��AfC���ŉ�(ՃAQ�G�B���\���m<��P��H��Mof+D%/u�R�}����"�R��i�ۘ���AO<_s���)T�ɭV�3wPk�;Y��P r}��p�����T��Z�W�u��Ọ��آ���[�7�*�Y�ee��_���p��_�y��u,(�\REٺ����Ɗ�c�|z��1��A�2!l� ���g8��k�ݿ@h`��3�!|��r$�P��w��:=v)��oŵ���Þ��Jjρ`\���sjK��`j��Oz'�*����R� B!h
���iW+Ϸ�������s)��A �9,k�lٕO0?AH�����e���7��s�ϛ<����v�zY���]���\4a t���<`�����ϯ�?���r2�i���Sqaö�^��O0��H[� -�;I�/9��=S�IZF��+x��9���#9�@J������@��m�K����g����W^$����Nj-j�E���nE���v5P3a�So��⧧O~���o��8��Ǩ���V����W(��fI�|����w�����n�X.u���?r��~�'?�<�y:>�f�aq��Q� z"�M)w�i)�+`�bX�fX�_!6�30j�ɂT�-%�9�l���@sc��w�7��k���&�GF��Ӌ�rd��{E�E��ܺ!���V�)0��d�+�n��]V{��o�>�lV����iE��>E����xs��HD��n�G�NGT-U`�%�W��,�z瑉����9z�\<RV(Gi��p,;���f��'����������\F��-��^�U#��ĸ����T�ݖ��� �BM1/۳�����@�j��t�˹�L���~W�-5�v��t��X�`�f�(K0�������5��^$`�4Y�E!F���K	����hg@aW�z�(�4��RL��0M�-��`
�B.tN�u�`�t���V��//��8'�3Bu�>�i�n�P	B����񂿍E��H2����vZ㇨8�j���I�LAQS8a�O?ˇxy[?��]�/l��
�$�<���;��1;6"k�G������'(_V3.�;7�#ò�ֱ�����e!�(�q3�[K;Q���r�$�^�8;�~�{ޕ5
/�r�«����G��#�bKU�P�P��݅����A*&uq7��&߻?����Ro�[8E�+-��lp�-�������ߗ��hDH.L�������	��É�*��霮'T5X�_�T��\��T�-uJ��Mfq�z��{%��b�0�.')L���X0	VFv�/�i%�'"L����%�T�8���69v�^4�4L
x{���sE~��0�?��<v����65������j���n�����q�#� �@n=�E�M��n�N�;!��1��mx���yL*=yZv����yE�w���V�~)k0b�ؖ��ћaTX�� ��/E�d�U|-fBAO+Q�ozfc���n^�TR2�� P�h��*U��$Im��|�sҕI"�^nWL���m?z��>xX�������� ��N�"�L���)iC�����@(�%J���(�`fR�̨��oظ	ң~wg�v�;�RT&��<\ﾱA��ӥ/$�K�P� XGU{4����r��!�.j,�������|
���&���.+O����s���v�m��Pŗ�a�Ȏ�4OTS����s��	����<�`Z���Nh5���T)�a�D�Ûl2�3�ݕ�
�(/bH��l��bfu(w��y? -OK������b@f��9�g���L�AN;u�.>I�h�%���Q \`���D���!Y�?	x#��x7������eStv��8{9 �s�5������V�ZK��w"T~�M�p��n�����D@#($������6O�g2�Yx����	OE���M��Y
���<F��3p���$u~h��ٓ�������ܥh�r^\$��%x�,}H�u���	J����J��/��3N�,j�����0��}���uI�?��
�x�y��=�������u;ld\5����Zɖu+� ���󆵾��1Td�H�I�hXUZE�5M�l"2��q�ګ��秕�}�llPa}¿.R�_�k+��h���Ei�2��Q�*�gyv�YN��a�������?N*4}+�B�v�I��(W���P*CR��ak<z��<��C;l|���3�����¿a��ʺ�c7��2��o�N�H?>�M��x�U�	�+���Q/�X�|4bb`h2ͧzb�9���[$"�A��"5�����UF@>0�����\�:�~S�:{C�#Xq�ओ-��R���ݽ~��9[B�������l#G�e5<^�K�Kq��3�z<�բ���	�����ԁr�x8��P��Ф~xN�O�pK_��ԭ�.m�M'I�;�xc�Z�	s����'�s?�ٗʡ�Q�0�"*�-7��u��h)�O�9���R��v�l6@��7<�I���J���H���b�����5�2~�b�T��7��Ȟ�k	����X9����FH=�����d7j�T/3E�v�*@TT6�Cό�q/��evݯ�'2�e�ϳ�6f��t?�r����T`2@��c�Č,[[]%�8�d�Q�x�^3�4!��'��<�Q��bK�|W�ȯe�TUWiFR5�s�7�0�ZjVU��i9n"�}����P�0��\�g�9j�Q
����d^F���3hH��U���������\������ǙlԮ3Ѐ�\K�$�e��h{���}{��UR͉���M��޶�I�W8��E���j����PFR��Xy�ix���It٦���C�o�n��e�_�=*Ƨw�[sz��7]n�p�}�)M��O�����#��$���* ��Y�CJc;bN��5�s�Z����,�ӣf�~p.��O8��Y�@.*������z�1��LWɻ�T��Cgz����]��h�)x�9:�'@���Ѡtf���J��d?�*��¤/F�t̂�����$����*���B��}N�k@h�-j�����ܓu&�ãy�9�)~�]e'�qm�\�����pICbO����<Ɉv��V�����aK~�������^ч��^)	g�C깇�"�wﮊ��Kk<�"m��QC�l4})�[�k'j&��{D����HmvD;ы�:IE`*�]�O������<�r�Ϊ'��l����^�����L�2Q�� e�|�~w["�i�Z>�'P�o/R�f���3�M�[z��.�&6�Y����c?Z	��J�s:c�R�t�T_p�$ĕ�w���i����յ�U3D����)������߃}�����0��qYԘ���q�N<uWﻄY�2�Ͳ���$5�g�1�ݏ�V.�eq�=���{�3�:�L>i���8gύ8}��Y*۾Q��V�O"��kz2қ!bK2w���-9e��s5޹8ǡV�2�l�Ggu2�}�E#�t��2p��X�~P��iO�w��x����8�e�碰"��GR� 6N,�0.p6�(lȦ��5�����(�0P��
h�����5��w�����Ǵ��ڨ��(y�� �b��Ƣ�_���u�Ƕ�^�]F��	s K����Ϟ�� ���]�8-�!`��4i�7%gR�z�c��E38!����,Т�����n��]����,S϶)~��\�{��X\Ԟ�1���2��ֵ��]�����6��/z	x��AvOB�&�y�a�3�9ʆ��G��,�p�����������H��
r'���������p����{�u� �N��/�ԣ���u�: ��k�0�y���zx�(մW��!�Z�.�66_yqAy��s6:���n�����<w7]󩂌�z�@x��n�6�U4����k�4*�}b�*��@�d�ag*+��ɑ�gTz�W�P�@!Q�#V���I5|y�!�?���S���12P/�Jg���Ru�6m6��S�`�w�g������ng�n��� ��B�J�Y�z��U?����O)j(���f�?(g��L��u��[\�iM=�y�!��3UU��a� 8����W���G|ܴx��� Ư�9�B��t���Y����_���P�lu��uk7�ԕR6��Xǜ��[����3|:��^�|�a7SV��_��Tɚ%�*��S[��>��yOKp�M7��Zl���J���^�;R�/�F�Z���-gc���NJ^?D҄[��zy����H�e�Dd�8/�qqU�W���6�OsӼC	�;p*9�vyp#��X������,&"�cH�J��i�[:�����
��	ô�/�1t�`��� ��%��"�.'�л�FB��"|�抿d�u��F�Wd[v\\W88�8�n��բAzE�J+�Hic��}�搵�Ŷ��~�;�?
D���9�fP�J�@���~��WC@G��2�q��}?Y�Ϳ]#|t�=J�)�O�c�g�=։U�y�̡%ߥ�sĨ$j��.��:��n0a��[0Mv���Jp��3&m����wG�KR`JS��&���.y�/th���R�Y���΍Dx��i�)�B���V=�]���/����G=d���Z{[�At1N[6��ՙ��#v3��i��X��C���� ��LfV%-#�C�����ڿy �ؽ��C��[��ަ{���O^���h�g� R�">;6j
6���6J�s;��c}tv�p7!m�9�qm��c�~`�N��J/)6�y;?��
�_���i�|D�'�o�N-i2���`�^�)�w!�I��Y@�,K����a r�T�&����5`�A���U ���ⴟ�����M\�n�?�g�%��!��!Q����,�w6ƲB�x�ug�5A����;��,)͵P�FF3��>r��璘��bj2��������q�l.����/�O�+�-|�:�p`�S��le�O���u�qg��f�����lV_�����QXP�Y���ʳ��l\u�l�Dk�@)�2A@,�$p�Ў�i/��P����þ�S1)/�T�-r�tA0���,�����:@��2y . �4�r�E'ڪ�o\��h�����t�n�&[&�xF�V8�j.�9��v�V��]!�";�vyg]����&�鄂E��
2�97�����z$鋶	5�*��[��bt��ա���a�c`}�7�U����*�X�tAjS_3w�.�)�&�]qw!��(���zΤ�~߭8>���nsg��X���MtK`�M4��y3i+����;9�t�|�#[� V���Ian�+;Iɤ�lY^9�qOf]�0@� f[R��7�����E���kK�C�/n�����g*,~���W���^6`s��<�/�����wu�ڬ��b�!�nhx){N|���0J��l�­xL�8�j"��\��Q���.�$
�y�D�
r%�!o͹wɌ6�H%� q�f*t	�j�S�L���I
*�H�b���&dz�ܯ�Ʉ�9�7�B�|�0�aq����~�D�U�F����I�af�� y� �O-Xs�H[�Y������:�i�q��@'𿨜z�kUU^�)����\.Y7研�fzs��]���\�{���I���˘��I�j*�9��N\�Ѧ�I4e�de���+�C��\��᣸���s�=�9=��j���K�@�F��eE)�(MKe�[��o�(ju��\��C�S=��2�l�G�j���6+i��&:�K@��6�/Ul���8-�kJs�V�ԖYrU!����S���By���]!�N;���`JOŽ����&�
�L�R�AK�-�m�d%5�<gl�h0�?�Ђ�~����i,4"ڭ�$�*�w!����-2�>��q�^`��p��_�`CS1wO�-<ȃ��>�1P+s�q����M��'��>����Ԝ��X��Un_�1Ј�N�BV�����S�vh���>�2�"49C�`����SA�A�u���0�D}�H�Wl�� {���Hv;�J��~��'V�x���
VM^�X#a��hds��:���ŀ�5r�A�W-.@��1S�/shy�2��6����Q�~�aɆ2�������)��Q����/��l���$�%�2�~��l{R�ٟ����;�7kZ7 ���֯][`�d�L���ܰx�v�^�li�|~����4�~�o<���q���A�i؍S��,`���������ŨFzǎE&^Z��=��<]���
��BY@���n�!vun΄����E�9Dv�g�{��蓮�MZ)B��)�⑼���6�։u��Rg� �����;��ۑ�3��c�l���y�~�Ye�����n`��T��_J�С�|�h�� <��7M�� HXm�5$?p��}�$	ˠ��FI7ӚR���V���=�����E������;f��,�nq�
x�b��Mۧ�l�P[T�p�A�*$+)oQ���@�:���O���05�E�ϣS�ͪ 3�|C�rH8ؠa�	���v����K�6�+��V�tnU��� ��.�TKe�楄�=�5r�O�~>�#wF����`����o���p�q�	�&⍌4�*�_�W�l���%	���ze��t�����G�$�\��QŲ���}��bD��~2nΧ��۶�W]��~z�4�x�9���Hk�"|v�-ש���\��Wnן����K!G�%g�ک�f�Z��[9r�An�7�%_A	��F�������!�L7���qmq�=a �H�az��p.��I:ܛ�3�Ѐ�?�M�
�L�1��|�kt��QU})kM�P�?��L��Q���W���9��hU��Ukd�+�~��a�pP�>	 ʪb9�^<n�3b�la�A^d�&t'��p��e���>����;O A0Xϰ�s��A|���-��c�pC�[k�y/�~IUEt�[g���l�D9��Q�mEz����bN�}@4lQ�K�a_�!%;��/�[��ƊL�D&�%1�T�����9D#K�Q��,��Wk�-�(2,=��b��?���YV�V]F���� �-�[�}@�X��^��+�J\=�r��z��ݩ�������%Ê�R<}|2�G���<S��ޯ�O?Y%��7? -Di�Zl'̛I�4ӊ�͌C�ױ�K��Q�V�k���@�+�}ٽ*#�st� ��o�����\y��tg&D_�_"qwv�	���]񐟳�z�-S&�,�	dZAˆ���~X��xV��I�-('t�PR9���pc���'Z�1i�ι������ǟ\we� �����+{�W+p�m¬�_�+h�2�*�(:7{�ɉҞ�*��|������@؋���>fc�v\l(kA�1�+ŋ�c� i0�oy��\@�"�Ú�xŪ2�x&�;L�����a�N�p�M>Z�֪|��*��Y3�9�k	���^q|H$>��Ö0��	����=7`�\M���Mؠ�9������h�R��כ�l��_U���s;>F�ס}�F0��e[ 	���v��C0nɦ�����1&�v ?�`�F�Iٕ�hk||���k��yM;�����}��?�7�����ƥŇ�dl#;~1z��8.p8U0N0`@ȧ.�$�2�E��p�`|3s��u3_>M�I��4u�"CVh�g\F
H�#��޶%�v�b�@�����H3�Z�$��~	:�5�J|�|N�*G j&��ɤ`Kr�fidt��:=����^V��)��/6�@��a���p����!
�Yn��3�j5s��\߯�")��
sM7p���B��4�0�>�����nYH��99����H���.�P���=��E�[�P���q�\�}�����u�'���AjqMt�����aV�s��0�D�@@K�s�����B"U���-"��uFy�x���s<I]~����9Ds�&g�}��q=&#-�x}�DN������1%�Ea��I���#�2���/��YU�U�+b~��/>RQ���i�'�wS�b��ՙ==G�����W 6�R�dM��c�����\�.؞jd�4ש�J䵦���p��߲1V��T��o�@�^�.��F}�j���8�ì��p��,#?\���c�߀)��? 8�tc3������E)��5�Ռ�?y��CE�K��;�˼d[���ePo0����1����`~����M��*5�Ҋ��U���)p�y��������aYz��w��C�s�ͻ���~c�Jjd�+��Xr�PDj���!�f����!�4,gi�o��~�oբ��-�}y}&�x��G;f����9��F}�6%���I45��n-�<�[�
S�I�xyMj0�B��m� $u0�^P�%5��YP�Y:����O�]��u�G�7���֎J�3���	�~J��?���2���V����~~A,y����Dui*z�P�X�������;���H<�^.J�ٝM���{���0Rt��_6���8�?`�wܖoFc:��{y�*�[�[�.��#a�Fd��� �ˤ˖��6��˘����v6��Ɂ�VX�J<��(�*�*Z
���K�D����r�C�(��ʄ$3�Fy�m���t�FGx����7JA�ă8-Q�3��I��F��&~x�g�~.� �ԩ���5T�@�2�Ot�*��N'�\�k��	#PIb��"�~UՑ��949 Oa�_���U�h\q	?(�F�$a�3�%��.:����Ob�b�� �Tc��*��i0��2��}� ��9F��xk%����8�jR"��N��:S9��f^���ĩ��������������Z�^f�������t��Z�Q��ۥ
۔���wXF_nX����eB�C���u�)��9�?I�($���市JIZ�*���
��q�K�P�-��e6@�JH�~��b�iƖ73�ËS'3�ɭul����EV�-�
2a��OMKݕ�$��9�v�j���G�|����˨�k�:`��.��o�����YVtm����D��t.��y��ȩ����[u�yK8��А�e��r��VM_<����:�%��	���Q�_qĎ%�m`�K)R[\r^�Hu��	����M��exm
w�o��X��B���<� ��6Z)������+,w�0���sL���6����[X��$j0�0�^���\����c�mu����q�P��0ޘ`�3A� ��C�[Z�1�q.��<T�y��Kn�m�)��nK�&�{���3�:
���OS�s-�ى&��,w3k���������x�u��ȕXFoK|������ӿ�C�S饼/:�|s-��W�(&;(\iK��Zl��-��Y]X�V��Zdԇ�j�%kZV����M_����C��8\�+�9�
a�!;�^����R��6$�g\�v�Ϗ7M�f�]]u��.��-��2��0�Ж��Ef���9u��?�v�Ĵ����=E��3&+z���!M���8r�&�ZJy�?kb���=
���]M�cN5~���q1̧�p�\��~���l�v�FZM̍M	o|�z��X:�ҖJg6�`�F����c�o��Jh|L0J;��jO<
ZT��5ϥP4�h;�Y�b�����Ƙ���z�?��ցXBY�)�U����P5q���}��hz�,$�d�p�9�2������[a�楉r^�f��2��1t���H��g�i@hPW9fWc�4��1foGBLM/��G�>�J����V�TymO�P&�Kv�	���`���}���}�\��L�]�r��=v�q<<4L��@�8ʽM~����sh����	ٿ?y��e�R'~<'�-��B�R���!�]3N�j>'����c����i����x�4w�����6��7lN㢉F��y#w���F����0<���o�Q=�k��.g����8O��y���i�1t�ZZ��؄B���֜�/2����=w!����l���[P��T�4�THt�N�Y&+�]Z��y1���C7bi����U.nx�E�pZ���(!��}P��0����^_$�6V�
��� چL��~Wӣ�O�2� ln�F%�X�����/�gi��������GK����I�'_o�>@�q~Ϻ o(�G�������h�Ak�ڊJ{�)� xM1�*L��J�E�I�������	*�AY�Z2�B��tys�H�̶�����J1T��{��g�9��.b������18f1Y�}�������l���+g�s������oC �`�\��g�(Ik���9Y@��r��Ɇ6� .����fA�W��L/�-C|�Ƽ�zW��u>S���%;Ɗ�"v<�fr#>��5pGnu1|�������2��a"=��B�(�ƾ�9��
y��鲶�\˩·�J�\�8 _S�pL)�y�A|�)	5.}���lf����U�3�{*�i���`�Yݎw�x�V��U1�5/����%����1��c���W�b
�����+q	|��:6k7�����1��?n�D��EI]!M�N�l1�����*L�7:n�5,*ɗ3�*���n�6���+L����U�n<{� |�zn[UW�#q��M�T�c��Z|�?����n��Y�j��7�y����)6/.����IŲ�����}}���x�#;5�y�Ai�#�
kyh�=�]�I�#�;={m�2a)೏��I��̯2�����.�p����^CI*׃o�Jw`E<ؔP�Y�NE���=]�0D�LᏍf��^Q�`=8!�ā�YK	���V
P%�֕�mV�4�
�wa��T�~� B	���m�1Wd�E�>���|�b3x�i���z��I'�����ld�˱"�CVʐfB�ѻ�&�!�4T�����sC��������}���}h�
ˑ�P���N`#���?g������pl�:? �v��4�yN��M�ߕH*V����?i#2�,W����gم�)���kGh9kO�T��Ї���\�z���#ʒ�~���r������%���f�	������.��n�"k��^�ż��=-&�2R������B���Y��@*��0��C)9��Y@t*��Tͱ0����y��}W���݊�Ʋ�<��} 2(ztz#6Uً?����p�A�kG�
"���>���᠂G�̟���Ǖ"����*�!lЂ��,�j,M��;Q(u�?v�j�N�z��2D6�>)�Ơ�9��e	�B��ä�����Y�	|��y�
SA�(PI.N.!=�s�X�yp�R+������� q�`��.].Y�؞�*��l�z�fyx�7��>�O�IY�����p��E�%<��m}�^"ܼY;���e�o��,���OR�Ĳ��aX	`��=���yv�aQ+sv$��L��v�ӶC'��ɼ�Ԏ��8Y�κ���^���L�ݫ[ YR��>����b�!.\��~��O&���#}md:a-"�~N]�H��-@#���6`�8>+�op������:�y�L{�%�	�:n�Ŏ�W	��y��C�"���Ueq��=e��D*E�E9���5�̤_��4�ښo#�j��T�g�P�{�Vd|�k ��c�4�_�g�7��>���uk�HW��e�$E������w��=�V�$A�҇���|�h���R��f��^�es�������\SJ�Xͳb�u.�Pb�B,�ه�A��c����E*@�,�;�DG�_����ְ��iWY�h�����93e�F���Z4��vm���͌	A��9��P�H�H�{&F� �XoV�?Wb3�f�vA���ѥ����������X�A_��N���s4�(�'��M��8EpÝ�>KѼ���bvn����)]0�4�\��jUd�l�q)c�W�T���-b�� �^D#�����ǟ��s���ۭ�=��>�Hފ󢸌�fr�80�ܚ
��UʊWQp�����":�d/�@u�ɿ>��M�(�+���1�7��9�ez;���N���ٮ�� q�%��B��/ʌuǣ�@`˻�����(���մ~�х٬��x�������3Ik\8AC��ɥ&��E��M<��,ɒ�/��c�;�:c����v��S���[���z���KHQ�{:V�>�[�� ����/:=^�{���z��nt��^��|z�ݳ����W���%�n���DC���)�?�cANS�ۤWG���m�$ۊD��|���~�1ز�Tjn�� AW�Yb�q��І�s�&�6CIJ�z����VU�\`E�v�>xN8��5pX �H�_���E�/~�����te�2�R.ӌ���dڙȰ4����GUra�@(ӑP�
�l@ͺ�&�Ƅ5g1�-Br�S�Δ����g|���M��mX���������.y2�Z�J�uj$�4A! ���Mt5a��.��ë^	���笆������q�6�76I<�[�D�^K�ҾTW�E��i�<x�#��Ҫ_�w�r��I�r��e��i;�	)�@��\h�g��OM�L҃�7z�W\d�ź�y���@_�,�Z���-mBuV�$��#SɊ�0�]�d	:X�G�x��	���M/Û����9��A���$�ȡ׫���J�yڰ���k><F\y�x.�n�$�?��Z*��4���]����N�Iz�G�ٸdݺ��qn�8)�_"�=/\�(Q�7�5j*a�?Qw�&m���3�8L)�u �E���a0kܓ�_�N*^5^V,@K�-x���Y�X�Jc�H����k��~�>����.�{���Û���KS*F�{��3�`���5G�Gk=M�"0�Q�lc�>��{p�Yc���kW�O�#�ڎL"_����k5��v;�+,�db� ����j��E2�I��g��}j���z�����������aryb�1���ز�%�W��:�&��yq�{t�,ޔ�4�o��7|�)G�+WYv�����������%�q9��j"%�Q�FD�k�#a�nw�S��c%�<�s�.�σ������HK*��
��ۺ���4��0���.g&����]�����`T�MC,z#!.U���:�r2�9�D]��U�����_��6�Y,Q�Խ-����!4�4�["C�1Lb5�"ھE�֢���S^�\l�85$ٴJo~Jw�X� ��ʹ�Ћ�L�z�DN �÷�s��^�����h0Z"�J%�A�A�O�iI��Tu!O3ǀ�
���Z�8z;�H��i�XEr�xm�����%�(A��(�t�ϧ=W��`�����=*ŕ%ǏU��ӌ �oM1d���^w� �*���Y����r����۳I� 'g�`���Fn��̓x菸��P�x�'�\c�Wi��tTƎ�u��=�y�,�]��\)���xk���\l*&�e����C����O-���Z���O����#Տ��q�=V���y6�Aoi>��4fs7=����ɸ�U:�'n �絎{_	��#* �h�$��������m<9���M�Bi��w���	C�,��E�k/�u��.�Qj1����3diĸ�9����!�T�<�l?B�RV����Yy
��qTx�c�����d-�9/T���K*��߹Ɍ��}��kd�(��\�=]�L�+B���E#���0�[T��YmxI����:�a��`�^};�`�F҉���CH�a���D�����H�p�lD֦�ҙ�8'��M��p��u�5$�G����Qp���9VT_��</�����﾿K�_گL�=�4Ǆq҂���1��)s�J3��J���r��>\f�1V��X�ܭ�)��&���'��D�e�6��A4]:�"�;���6��4�.��E ��r�1	$XI�I1���{��.�_�yuB����i]nQ��17�V�q���mю�w>fض,�	��j��NS+��
���w9\>�0�r:��T��%����u���+�␼�k'@ź��i�n(�����}��[�'{��X��#4��bx΀�t�V��Z��::������00�������j�^��(w�t<jrr�
oK!����ѱEw�f:��r=
���6xF#�D|�z/�����=�4j��~bF�4����mCj�CT�^�z��=�lp�˥��abC�"1j��{�'�.�7m��E��\dχJ}#e!�_5V(�E��G<�<�X����B�hF�?� �͉���[mu�����|�u�N��uK��y)r�ز��k�$Dd�ճ��Ñ��jF�����F���ud�D�����T�kx�W8&RR��d�%iCه���d�/���%u:!�b�J���P�Z�����W� :O�~�)1+
@ �Xc�r�9��$"�
��ʲ�q�6�Lm��|�0�M�q}�N�3E���%�];��#P��3�p�k[���Y�>>'m�;�^���kW���������+� �x�ji����u��M����[M�XR<�����B��be���-pٍ��L�V����S�7B���hK�w�~��c#��e����S�
tmxZҷ�0��C�aSqL���6�0��D#��h���m!���N�1�
SqEZ��7�D�YQ�����fݸ�d��ق�]��5\)���pB�
�QEb�2��/9�<run�	���T���h������s����p�r�.0.U�I����}�i��n��*kia�S��5t��|XXYqR�e�29P�ʭI[��,Դ@��V�FZ�ZD�~q�I�عUa��|�ɈZ�M�4�k�GO#�
�d+=��cŕ��9p���A�>�蠍)�Q�84c]�������ly�5'R��e�M��Y�1�y[6������@U��3)�X_����$��Z��70f�V[]�9���Q\��l�8Z�'�����ۣ��S�7Cw�.�D%S��X�+�?al�H��x�洧�x�ӧ�!�pUi�1³��u��ܲ-�?!�*�`n>����T�)A�2ڰ;ibi��6�R�3ħ�������©��#G��4����}�r����>�4}�XT��`}����'����nj�茞�`O���<�0��ڹ����]S#c3��Ob���{�Ќ��?�5%='�v[�M��O��`]�����L>�y�n�� ��-������͍�!9<���l�괇f:	>�N�����6s`� *�MTt��14���_���j�sP���8����w�I���媸�s�膇�dg�3�<)���^�v��Y�5V1�����o��F�a��Ø�{_Z�=��c�2ZG�|�]d��]xr�5K9�ހ8f0�8eds/4�w��dy��7�qj� �g�G"hʉ�OlJAO�&���:� u��z����H��[��#��od��zX� �4w�늢���Um��Z���]1��1'�]0`-�I*~��U����T��?Uw0}p3�up�*�8	_¬�`���@� ���r��+�Mic|#�/~FH:|��t$���3I^��� �#���ľba�xw�Z��r-p3]�y�uF�j��*#bj�S���&3n�b�D}�@d~&\�KX��;��B�Uo	g^g�+	6�Cm�宲�'��߉;,��^e����aK웬�Rn������2"�#�5�Z)z/�Mg&��-A����QT�Bk& ������H]��+��;t�Ǻ`⁤�<N�/ZAs��&���\�K�Df7*�g���?qaq�����-��z9�����"�g���4=~�$�w�\���Q����C*��o��1��X�P��ژ��iz��y�53O�,h�UX[�"?%[�Af;h�)!7|��}�Gs*�zT	�j-�;�֔@�d3�@.��5Vko�K����'�K��%\�z���i��
�\O(<x-+��[u|�u	��w�Nk���\�-��8"V��n3΃��ie�g{ �x�(���g��j&ؖ�&m}���#?�<<���0�'G2��rБ�PiHa�
�{��2A������
�R��?�W8J+�#���Aq>�H�I<� h,Z8�8y?��A�9����p T~��*R��cWE��!�q��(0���9>�+�����vA�����j~J�R���I��cb�T�߼�]���ZOJm��Ds1Ҁy�/υ��z���c��4���P-���J9 ]�4�ɟ0wxm;��͠b璮\_$���Ž���%������H�'육�������������<��uՁ>l32:qFOH,�1ʉ4����F8���c&�AJI�]�g���/.�X��Z�JGG*n>%���,�s�zCQ��h��!.�L������z����j��(1O������kؐ�K��Å���--v��7�i����+�U���z�D\�"����\�:*��&Pj�n/s�'�:�Z�	L��� ��q����~�3�n�d�g��X>��Up��D�+mW2��[�nU��B�q�V�wH��/�?��o6�]��Rr�,#�,̖�F����6�O��^7�B�P�(�k��/���U�B���]��ez�K���YX1�&"P	)�8 ��JsF\ 4�콎�8#�=�7YI<
�4@H8L�0-o)qai2��x�
,�2�0.dF=������D[�N�6/�0�[� �����d�����yUSnD�ۇt��V
~ 	b�o�'%><xw���F�u<�R���ߜ6.�z7w��8h��In�Ə�֕x�zҖ����|Q��U�ь���5�
�S�D�LȽ�L�ou����u.��-�+�"�ҰڙG��e�8Z�����m�%(tp�=�^���K�����`��̠mv
X8�M�1��5���PJ*��氮k�Z��l�J����i�\����~k��\!˧�H�[��u�
 :���c�J�%�v�-1p�U�p�n'*��@ev��ET�cԗ�3���(�(�8*$����b�Uj�M���*�)w0k�XsxCt�"��>U6��x	m>/Gj0Ak�:�(1�j�E�U{a.��P����~��`8���:>�߆@�����D�|N�XK��[H�4�#�G���E/���>`_��t1�\*�#H�����uS��b~���	�H�*��"��5��������
�$�9#�0v� 2efA��%�&C�cB�1��u�wa$p�T�Cp�<��t�9�==3�p� D�&�ك�{�n'�R<���ȏpI����<D���q��B�N)(Ά��v>��y3��oSv^��g놿Ԓ�_�J~ �����;jA�ԎS_j���2[G���s�h�vz������5��.�]���3�U���X�cnx��-���i�1-���V�<O�k��{`�+��Jd:�f��BEb�=�ɲ�T�F�
�<تbW<�m���m0)=���_�$�-^{@TNV�G�� ��B�?���}Z^�z�Bg@N�ϯ�Y�I��_m6����hB��P��iY�5W��h�� Z5���S�2tP�-m�<[+��W{� !-?O�1cl���ý��}x<FV��4u1�/��?�;H�.scT7��0X����Q�8Ԕ����k3d�d��&�2�Ǥ8��w���C�va^�=�.�C&OQAE��n���ejw��S�m��Zrj�u�\ۗ���4����0�|�i9-��
6X���l�Z��=� YN�z0�	_"��vE���a�2��f�=�e����$L1HĦ�TK�CQ��ǽ_��(��[�Xii�]�j'����h$�y'f��B	��ٿR+��@ű��,�8�s�����(���m���H�����6�F3h
��s�b��,u��z��"�$�NX �h9��W�Đ�*�y�|p{u"�9��z��d�m^�a��B�5uZK/�Z�,'c)`h�
1u��տ0��|��`��=�~��t�L��_s�5��� ��Y>�|v?u�<kUHd���H��`fu4��t7V�S����Y�u�ߕu2 5Z]�xj%V��I�YL�ĳ�f*|2��И�(֕��A̩�T�qo=�����$]x��	"d���T��g�Xq{B���V�� z.����>肺	6�fտ(�U�s�r�ត�*#��G��h>�e=���a(PR�M����rN�OY� �ݹ.x}�a���F�%��y7R�'ϡg��@���H�6լ�L��"��kO�ߨ@V�B�B��(Ği�Sq'Pr�#��tP�2-λ��q(���d�r�:|��M�U�}I "�H�틀C�ͤ��,�r�ͣ��fe��=2�������\B�;�޴���?OM7ϧ�L�଩�̸1~���2�+T=�V9<��!p~�������r[ÖNT̄2�v)�RD���N?E�j8��:�+y)K/�����B�V�hf|w!��f��e[�Y�W���]'rε��ە�<��l�������)vNn�o^�|�~
͌��w�N�w;��$�2�0{�¾E���[��Ε�E�K�A4R���cp��i.]n+�e�s��7xU��s�Vh��ݵ�o z��:�*(�����lϽ��=�u��έ�	�8O���w���>�4g\�XN¸>�S`%ʟ�R��|=��~Ւ�5Y����?�.p_U�y�7-�5���Q�F��$���U���~��4�R����+l�j���d)����^WL�P��a!����Qj�h������:Vg�D_�̍���������TH�ߡ��FpS�Cb��:�p�"����ي��%oO��dn+K�`��\���vt$,���SG����2��Y�J�C��#�ϾX<=��Ó��|O�f�A3�f�Rm�}H�
{L#�֟�[���Yĺ2_�հ�g?ˠ8N�b�4_�Z0�T���r�FΏ��>K�&��������˩Q}kR�<��$72v���\B����sNy~��	�FS��㙣�}Y��Vm�-B�TO�f�t�N�]���`�4��'������t��N�6n�ꧠg18L���}����L���of�a/��Q��}O��prgg��V%
L'*������~�E���-��:��%�o��@\M2}Az��۪������ @�Q%��	�`��/�����1�!d���&�կ
��,
�؀׃��)_��?s�d>������wBe�۪����r�H�D��f�%�6��'�k�!w!�2u��B��E>tM�~2ft�+6<+k�S'������M�2�<7`�loCy���[�Ŵ�'	H�J�ޢs2+��^L��߂��A��^`=�Q�@o7��c'n�*��޽�o�`F&�p���!�����}T�SC<���mM��wM��5닻��P|�5��h� ��H��
Ǥ�����˾�C��C���e�w�06��>�>b�,�g+�zf��g�PNf���U��B�n	2�5o�̽w�%��j�k�Ů�H!�z�ް�T���3���:��W���-h5�ֶ	R����dJ���<UϏq"�eE�VV��q���h����.�ͪ���/��p�` �8<����\{Ƅ���z� ��*j��d���8�:�V�oh�6G�8����l�z(nc;f� U	����5�=�"�`,��̛q 0j&r�д�{�
*��I�AT�7�:���y3;%ir���g����EG����È�Nj�&��2P���ֵ��>2��@jZb;�|�]ӈ���/	w��I�BsuJ78�O�(��骵��ڷ�Ϝn��k�"w�JnY,�n����cyn��X�\�o�����e�<�./-_�W�f_�� Դ�m������~u�1	W�H5����́~8��+8�������o$�V2��r��~�)ߺ�Δ=!*m-b�!�ӓ����<v��	��X�2r�)�[0�-6��v+�~��'30�*�	�#{���=�y�?��"�RͰ��D�W��[��h����'��:z��zf��Q�Ou�_9K����� �L��$�>0+旚2�LF�BB
�1�gL��qՁ�
�뻹���Z��+^��eR��[�����+#hI���f��������}�N�gn9�q��,i�츹D{ ��N�"�_1�n�-�=��
����+֦��������
�T^<��ジ'�k��~�""(���Q�^v=C̒r�݊�����@;J�Ʌ9�G]�K�m_=���*�C�6`�烽i��oV��]�@���z�_���R�P;e�12-�<z�E
6T X�Ò�Τ�4ܨ�V&����W�xӹ��������� ���)�j�8&$�x=���7��o��L�F%�X~�كz�"T����n��J!�9ٓ��G?{�DwAJ�Ц>�%�	��}�����髮`����x�h�D�B�+7���i!��$	Qi��txd-�v߅��К�t��e�v��H����_�����O(-A�Y�/��y_b>�
l�����+���M��[Y��A-�T�tt����ZA�N�xFF�oPC��o�Ҝ�\@x�1q.�b�����=\���M��!�0-������S�Zi�k�"���GV��IGjz�{�@��0���ՠ��-��QY�^@@2��QwI��Y��?�\�d��i��m��y�۔ ��3Hڴ{���u�wp\���(�N�$��I+*����[ّ7�"2�z2��LF����G�o�E��p����eU��!�A�Òz�N�����zC ��V��,��*\���C�5�qsâ���f4�6�k�A��Q��P��Z ��?�-~��q�m*ाQ�Rn���y�P�cj��Fw��k�~��d�����E�!;3�R�i�����\m�����^��l+�O4g���8Vm&��`{�|J�m7������V�p���[�΅+zӶ��ʘ���@��~�s�"���yc�����\����;��C�Zli��]%���;����o������̞���2�>6�jP�I΍�	�p�%�7[��V퓷0�:����Qc��C�|^��I{$�P����KI4���,f�ܟC�^��0,6@�f�3�֧���銂k��,^�O��V����G2���1�oMeȴvmC��Z�O=oyS+��yBl�̈�8�ҕ���q�m2�dz�{���krmLwM�}`�d�<�-u�	^i�!�[�։{0��U}PR~���%���7*kҀ:�޵X��|E�*V���j�ǚItJ�*�(1�G5'[7�qtA��g ['�����I��?7HV�(�i-�\��s��BWa��r�.�k]��t҅&`��>�R�
'���,'ђ�܏��_��@z���ޢ�����K�z��xj�)>,�x�]WU����w���vF
u������,�M��LN�-�Xwq?�2=���@�����00����~#��ȟ����A)�^7{�L#{u:�c�u��SHR�<�Kn�-���nT��7�ָ[�D��sC��a�f�RjSU�>�M�""�%�P#��[A�}s��������(�5={MM��=<��h��-eYs�/�\�}l��k*�E�=!M+$�����-��]������D@7q,���}���@%�CX�d���(��V?yZl�1�o��m����8��X�"���x��o���E�����a�O�������)��,`��!U��E�"�^����(�W��.�w_o]�GI��^y��@֒��Q�O��)��^D���*�����p�Kɕ+j�IZ��1H^w����<MG�f�d���uu��O�zT��-?l�X"�ǉ~�եM�]������&��<�T��wD����V�_k�5m���`�;1���}����k��߸����E��J�V��±cd$R��T]��S|o���KiigR,�Kِzx_�p{����;�]!M���I�٧q��{��m%u!�j ��O�6�e�T�`V�n�f+�uE5�<:	�7wc���/�cM�e�`������
��}�����R#Ŗ��?����r�05D�S�U�;��t�=�%�]�5�4�]4�[c�Ò�T�-m�"�n^/^���z����A�$^)�w[��Ob�6��9X]gZ����tH�ޚnNJ0���||�k����jy_���hYT�?R�����k�.M6�C������{,��. =��v��)�v�9��Y�<��UQ��p˟�E�z��L��#F���3��"|O��;,���:b��{y!�I��gC��vӂ>4�N��Ae�;�����3�zk;��G	a�sZ�$��[]�L6�@}�m�!^B���h�Lm�K��g���_^4��!(+$�gb��|��A���*�ي��E*��;Ã�U�. ��n�aE���6��Jk�(��PO�wS@����-^�U���q�"���#FIj�4�@�IZ�?څdN��
J�cx6� ��c�����-������ ���_��
�\�ӫ�`q�"�O�<���t�a��ZͺZM�=�\`�![��
x��)ԁaDfW���/�����ۋ����J&�5}z�9URYn�J'-�mp�̎'r��_���7��uzu�����u�n������}m��~�Ǒ h���9Z�X��&i���~��T��n���w�P6yŸ�'[]���r 勬�!�����J s]y�I��aBÛu~��G;�DE��c9p@��Q��u����z?�߲�(]\dp_wk�͂@�Lgh��|��?7V�xp��%G $Fv�kµx1�Hۯh�ոG�sZ3�A�� 9�TI��U��dj�6|����[D�����}�LtII���_�*�z���q���q�|d�U��{h�5��n��|�\&�;�ϱ�Aw�J�-��m�B���$�wdE�!�;3M�։g>i���@p!�$12\��,JoZA<3LD��_�shq��%���� ��)��Ȟk���H�=�m�~jx7D��'
�6��x�?o0:��TC`43b���4�`�l�KE��pPYϝ��T��Ǎ�Yյ�&L�1z�PH[��<�r���/QpA��5}���>���^��|4x�-���n끤�ؒĦ$]R�g��[������>2QmR�*+�B�(�NeƘ��W��z��w�{Q[C�(8ʶ��?��L���e�N�V4�oŝhޙ�cJ>��Bu���d