��/  �-�߰B�P��ي�m���+8�KS�����B������+�rz���C�
c�_����b-�����<����.3%���'���jdM�����S����a���#�e	i{�E6RQB�^K�Ҧ����^P�~�>�=��zQ�Cn�OĎ0S��{c�Zf�BO�����U@G[l�Gݹ��W{���ȑ�����	e����Б�䷒5k,���*�'oP�'Fz�q�3�z���XۉERl�"�t�Eޠ��f+�yD�]�X0/���7��l��'��YŌ�=��1���^�9|�r�w�8�#gXN	��@����A�,��A�𞪐j�`XؾG8�S�F�䏬����tZ1I��Z�㓬�c�y}j� ��c~��K��k�\����n�-��[� ���4�"��B�=~����D��-�R���^Ƣ$����Y++�WL2t4?��>��=����,��.��Tt/]x���!;�\��[�x�e\6��،����ج8:۲ߊ�*.ѷ�E��\:Ϸ���1�x*�e�}��0�0��a�5L<���ݮ
r���\.q�6�����Ӝ������9����+�HEh�aE��l�O��:Xұ�U6n�Df ��y�J��� �ij�\�ΧU�א�)+)磳vzV��	�&�Lď�$�n�9@�:t:���O)g,K�[u��yΟ���0�A��;cV�IPK���U�T�L�8m���_�Ą#���U��Β,�뻷*@i��OϏ
H�ϯx�04��'�2Y�;e�g�0!�Б�O=��$�rW��`"�f|���J�"�j�c��놣#:*��F>��Px���ke�i-!��5�~.NԒV���IIy���dM�"��Ùg��E�0U<�1.V�:�?�a�f��߿��� ����@f#f��9q1B��z�s2kFψpo���c���:� u:�1� �Y4��[�(33�f�?"��EM�	�"��_�� �xG��O�v/H%�i](�\��4)��<6}V��>�Pq ��M�E���:�U��4�?��TDt��>��g���(�AV�$IJ�bH�l�2P�ģ�"�ַ��c�-[p�{2��0�2�Y�&_��+Ӟޅ��[>���VB�&���j�\�4x���ֳ��nS�נ�4qߓ�1�i���qjM����}�o��K�D꘏��B��|��E���
�g��t�{�m�T�/��,�����|��PF.DY�%S�p"�j��'��۸�̑�E���ٿ���Q�%�A]��K�w���N}�_0�����c�eQ�q_�W`������/	�@l�<��8t�Pg����)�{d��E�?o��Ϧ|#�$<�c�)c^�3%䠘�3b*�,R(��,��6ղ$���A�.���5�A�o,�ֻ�(o�Sm8I	
�0��F�������������(���1��ѭ�j3�1M�Ηq�Q��>l��E���Q%-`�#�d1�G�+�t����c�bdF*���4����G0S��1*�\-'5���6��l"��͇Z��N.�R� ���JS@"k0�M����`��K�R�3�EB�$�v�5rjZ�ؒv��/	0�7 �D�N��#c�q����A�,uT��ۧ ̈����&T��٧���h�}�
�o��¿n\MA�=kT,�m��0.h��HM�gK�S,�E�i�}��k��Y {�,��XE6)��)���� ��N�>nvK*�\֊>�,G|m�V�U�<�z-Aain��a��aCR^/z�F���K*F0 C��Fem��U~��S4�RQ=E)�M�%���:g�+q�8������0@���My<Zt����>�Uxw�Đ�{� ����]���b�Z���^�CQ9D�1~@��xF�f��ɔ�E���R]���Ayw�'���2��p׎��ʏ�T��KRp ��~��7/q�f�Yp��l��B�YK�?�߂]uN W�h��S�2{�Qg/��M�O�`POoU�s�/.=�3W��tC�^�ns�s]�,�eI>�4�;%�k�Κ�	�M�l�LE�50��WG�\�lޫ}GP�r�HqD���"f��byIo ��|������Ì��=j^�����"�K�W��IrM7}3#g�J�7�0�����.qz������҄�;2�a��i�#��6/�奟f�Z`#! Y�hu't����������4�'>R{��̚� ��xVh`�F%�!���k�?Qa�;x�w���IQ�������&A�m6�ho�V�����z�� �׭�Ż��^��?)m{ղ�`SCx{r��J�tF�P)>>Izw�P	`��ߧ<��(�J�Z���u;�G�d��m�i�zk���b�i.d{��f�PZ���dl���؛���X��$�'t �{a�)}��vL���g�T����n?T�^�����c�fa���!~x<��I	Ѿ�l+Qd���U�������F!3a+�4��*���E� F�Ů��\��j����3s1�
�նRB�u�B��|���4�o:��Q 0C�Y���a�<��¿:s9�pwȔ�g7ߒ6F���"�s;Ň�D���ݫ��_��]�ھ�Q��}��&3����g� �@̑�/����J�Б�Ʋ(�\^�E�qéC�υ����r,�X �usܕ��,*}��q]�3�W�A)�DeV�X��x����̙b���W���X��|2�~v�99+�!�����g���a��=���-S0Z�uglF�c�� W{�@���z6R�l�&���m<7覻o��s_N�Kp��}Պ8�&��i[2[i~�:;s<��L��tx��(�x�X�Gn��}n�ۺ[��W�.�8fQM��4PU�L�� ow�q�F�7_�Iqh](� >�D|�omרY�jo���L��.����.Y��ģ4Vv���ʱ}�֔P(�$f��z�>�|
!H�_9��l��݆��:Ub����`�"�]IGiT����x�:�r �%�K�0�0���p�5��-C�>t9�e@����(AvM[}Xp�V���b nc�����*��=�7J=�ĥo?'���/y��ͽ��Klw5��Uj}u���C3�"�����%�	��Mj\��<�n���k�j	��ڊ	8?O�p[
�ڐ�W��]����Kf�0���2۵vE¶�3��O12����-��.x)�ܳ����9�/�� �\�Ϻ艪�U�Æ��ӛ.)���7�E�$�t|�+��
��T��,�v��o2Tb4����t�?|Ҷ.���D�	)���Dj�Vd�u�v��>H���z�w��к����V2�G�ac�ຆ�����Ȕi:���Z�g�����f�f��\^?O���54q�s�B,�K�q������Κ 0�����)w>��k �wt��X>�>P��J�nJ�N/�n5����	�EF�����!Y���Q˕�	��z��֟f"����Su���s$S���]�e��vv�~�����uf�'���:`�͟�'��$��ѩc���'釔��q
V%
A�������*wU�pck툯7ˎ���i�qەʚ��o��<!jK��d�.�ܽ����=	|��l��x@��M����	�!֫����F3����ځ��)&5w���uJkF	��epnC���i~��h�C�^���`�g��C�5RK�:�!��c�<���ş�5x�P�@ص�-27�z���3"�G���BDƓ٬�LP�9��*��J�����4��hRL�NS�D���$��tz/���s]f�a���ĥ�;��^K�9V�-�ۦ����oN;j�(�eq��%p�#�ߵ���J��mR�ʶӠ�5^�I�3�w��\ {��ؖ����\�T�"IX�V�澛1��?��^�ff�jJP�z���'4p�T(��_kF�>K��M����1i<9.�Z:�)2©3�0�v#������6̜ �Hlr�<I*�A�4��	.x��W��nTߓW��"���v�e@����:��5S}��r�m�����<+��A�P9PnF$���E�F���0�F���]�p�<�- %������_Z������_�~�2R��g��Y���SFWJ�w��'��u?TRA�a��0�j�]���Prn��3�6'����I+�x�?��i�a�Yf�ކ�>�`��k6�4���Ę�9�/kWڝ\U���-*c7�t���d�r89�)��Ëfc��̓N����녖��1�U��j�|RɁD�dG����Z�ɇ_����������"�K4/��������?���K�ms٣��~h�����8��8�Wr¡!��,��Gm���V�ə��-��G�^(0|�fB*(q`�C(�v��~�f�lGv���Xr�7��*�C/���KC�*����^�	5|	lӬ���a��ë���@�M�-ɹ�J:���a&������]y�^�9����3�p+�x�?�����I;�E?�/��"-8+��I[����e��H�p���O&ۋF�����OAg�X	D)����,5����:M}�a���>84�W�U�`Kϱ��{�^�Fo��5�׏�,#l?T�1N˺@���6��K�'���s~��R8�uMPqF�Vy2���wƏ��t�@���z�M=�^Y�'IP�/[fio�����#���1}�;�S�)�xa��;�ă�p2#�~'��q�S,|({�|*_�nү����� :H�|u���G`���4�J����YΏ��@H�)|�P4��0��[�[}o���q;wb�#U�5�]d��k�n����0˸Kr2��C�*%����OBED����Մ��� 2Xؐrx���N���d�� ݨ%�as�R�V�Z�x(��W�*�@e�$��X��߮s�J$�j��͜����U�����H������B�����F(F��[�Ejdm vy�w=��;�w�g~p.��%�x_!� {��5{j[/�}�����./\��h����u�!�M���U-3T�����NZ�����8�e���m"CX;g����lS�����r��GF��w��=��:�$���I8U��~nڠ�*�˵-�qn����wg��f�VJ������ ��<���NW̽��]����yf�����(3�ވC�
M�?�ڰ���z�Lp�#8�t1h��7X�������<�2��,�`��a�ᅊ$"��rs���6��[���sN2��/�����E�eX�SM�v�������Wp�)d�А�Ջ��<�1���Fn+��5Ŧn��oR��^���b���ń�͔�q�M
�I��}��T� :D���r�O�t*��qUCCv�	�4���D�ů�Dxl������߼���X�|X�P|����l��o0O�\���K�����!�$;�h2���<�H�H̯���&��$u
] �|�0��4��c�� ձ���pA��z�}쪰�?/�RSezo��	Y���P�xs�u�n�.�b�+��e�����]վ�#ݓ 	d���4u%��W����y�:�Jm<��'�^�'����"��^M<Қ��z���g_�l^��3�,R]�dqA�O	��3u��-E�Ji�1�}s���^T[o�AvM���������Ml��su��N-
`�<oZa�Pj��D���G��1� �U���3�O�3 <��%�V��}�D~,Z�j�|���7�`F�)d���z��h;�c����@����S�n��?�k��ね!-!�]7(�����]�����!�ܖ6����YW}�f*َ�۽,�-��H	A��>Z����v���f����
*E�a��fؼ�G
��n��I��K���_�9&q*�E%����9�	GL�6{eH=�3�E��(�p�3|4���1=m���7�F_�C�"M�z�^L"��}�: ��0O���/ܱU���*���������!76���dڼ��؄�1��=ÉW�>ʀ�P����*z6�)���!������G���"Tr����v[���`��R��zk��ӱW^�H!x,.�n��yO�{�����F�������9RQ��,\ڦ[h����q4�7�b���O�M|ae��>��`���H/��˞aW�� ���i;�eHUι<��4��q�D�Ʀ��JƝ�?�V= �紾�*g=ܐ�/�����K�E`�]�<V��+��4eZ`���J�w0��8��2
__�vr��m��>�9Nl҉@m�G@`��x��?ú3�F�����k;m��g�v�x��$cc�YB?������;��5v�C�g�!A����;;5�+i@�,9��^��p�ծ!��qAB�3c�~U��E'���rT�^a.:����Hz��4v���f��r�,���z7�H'��M��`h���>�	&eh�·�D���z>G�?����b��R@f`i��l<���U��m�F��3�j%�\?�>����^�K� �}&a�q������#�sK�Q&2��6S��)��i&���-]��s�S�b���(� ���{����:Q�BK��0悜�n y�����t��B��bXr:)�}�c�y�!�|���b�䂿M|ѳ������'�n�^�j���r�t0z�ڜ~���C��ͥ�$�TP�7��B2�L��v��=�� B�g���Nj�_�X�ҧ,Į9p�Vq�:�v:>�yk Gİ�AX�ˤ-k�`��pY�|��q�Ɉ��iت���s�ЅC%ցoGJ�����'�^\I�c>H�)a-�#)	�ff��R����sA��i�A@ˬJ|o	��>.>�k���ξ��%ǚ��4�cf-��D���WU�~D��eq��������ҟ'n7Z��>CZ�ɾ���!	Γ�Ԣ�B}��B!��� YM�r/�{��(�r��"�_��R�-O�J�0pMm���ci�,��(v�7��½z�r=*�_ف�u���(ۮE<��x�H�"�1����Z����E��X�b}û^o0������U5d�B�q�c�L���6��=o�%�C9l���!�xZ(��}yf��ȝ`���6�6��"f��ZrQ\|��ϙIܥt����x{U�"*�wY�`*?i�?k��e< �57���3 ч5nʓkK�/���o:�W0�+�Y~T���)��|��X�Υ�"��KE,������f��=Q��Y䧫Z2G^��0�8�@����[>��M �|eW,2�j�}�>��*G����dr�f�ٕ�����_�i*�;Z�F)[y��M�vn6�s�7�ǀ�O��� �K�F�X_�=� n�.Pi���b�s|�
�ʪ5v�mh��'�2���S �~�����#������y�@6k��dܰ$����:!v]΋�W�L99���{X�$�U��a+�ͪ`2g0�D'/h��[�����?9�&�Ei�Cz3���|H=Fhωʸ��7�Y��M~=a��P�u�l�2����5x����P�!����*I�(�G�9)̗V�P��g��c����tǛ�t����Z:�wΊ+^3%fڥ}�΄�4u"s��1t��h?(w�q�j��C���y�������<I�2��h4��Lо��I4
��P���������n7e�Qױ�n�,n�$i�S�ҁ���f}���Ɵ��e���������[���1Z��(`LNK��uw�S}��&]��i��e;QR�(�*�)�
���qove?����f�<s*Ar��� D$|
j�I������pqÃxr�����?�]�[x�G�*Y)%�Uw���+Q���}�^bbf����C�fy*������0J�p�[CB\l��y\d���~�`����F7�.�fP��CSc�������0�j/�ҢzНzR���J��M��8��|R�7H�E�g����D�W��v!��Z�7ԍ��AA/_�0]�gDٕ�(�#V���7Bq�bN�v&TI{�4� ��I~m�i���\Î
�_N���[;�,�V���K�
�dh�׊[����9	���Bm�i�%uLA$Gפ�>8
��̏�l�S������ǔ��o��_8��<~W�S�a�J��-���l�:mņ�-�$L2������yŒ��jܣG��8�m�as��
������{�}�����r���̿�P��L�+I��'��E݈��Sj����s��VM.0�f`;{r��|��2$�s#���%Y$)���~������Oe�Q:�������Y��L.iS�آ'�W��)l�OH�H�|������C���N�C(b�76�˶��/��,Q1T������W�>=��y�p��+�~-}Q���'��+*�s�'{֍9�K��i��GjIl��$o�I�(ߋb�Z)Ҵ�_<��*4~��UQ ��:F]rij+��,��S�Q���Y��K���G����8\�SK���b:��1k����@#͵r��\ej��k{��F���.r� �H#��Ѥ�������^�����/U"Dn	ܥ�v��w����ʨ�����ާ��80O����Ü��a�iC�[����R�H��[��V������I����b`rl&j<��Wb
̄ӜE��5���s�G[���c!m���	0�����E�'��S#���k7E-�c���u���
�Ҥ(����P/���pe�m�{��~+ѯ�f�v����ń=�o����V�TU�̝�C�{���Z���,Rj�,�tjF��/m>�j����k˴��V�N*�Œ 8_��ё@��`���=^
�5"S`��6����|��8Z��LI��֗�W��Kv+S$p�t�-�Ch�Wk�S-o�LO����J��d�M�����ޙzLQקr�3��>x@
<M�������Rݢ,u@6S0~��Y@Ǻ��`��o>V��T-�������AJ�2`9D�8v]�*Q���K��;�-#JF�5%ds7��C�"�v� �m<Ruuo�߷}�2�ޖ�u�Pz ��o.����d>/ˠ�μ<@���K�<�d�7���nV������`M,��������bsʊbҡb�Y��[��'��!S3ʁu��5�9�穝W�-���L���4�<����!xjQ��`��^W?%'	�q4Q䔲?b�����G�BtFN���#h��sL�"}���t���r�Ի�����fK�C�L䟳@;h��� ��ƵTZ~K`����%�W8�Șm:~���Y�D̒5�_9��؂�e1����[�Q�kzؖ3����b�A�_��%@V�{1~��l�\��8��1w��b�!��[���X�H,�����ZW�Zu;�pY���c����Y
V�II�� �bnG��Y��2]
c7���+�.7U� �{(#R�HGA���Atlvע�υ�y.
�xK�Bt��°,ų�lB@Q�K��^x�N���
DQ�'��G��"8�)��RGy�St�x?M$Be�����cŞ#���k,ߠb����L��ξ�����6��ig���M��_��jxe)��v��&�)��xS�M��B�(��z,�w�.˂�^�<|Yl�:�fÔ���W�z�tT�;��&��nr �l%�(�,������sT�V��_9B�"��i�[�s�����m�"�% ��
�M3��͏�ǜ0$�ԭZ-�N��� a�J-���I��ȧ�Xdv����C ^��v*D >Kr8�_���E3�ll^���G��F�S�H����2�[��R��$-R����ijk�hx[�����8!f�Eu����lQϠ����e�rp�Y�o�?M�^��]k`�:J�ĚMj����s��f�#�S�+|��İ$e����ۺ�h`+��͌�|g<c�?n�-u*!�;15��b|��?7~g���]C��%}t�l`�]b+w��T���B*�����y��\�:Q�-�v�ᗎ۷ͳ��k@?�Ї���Jo	�-��xQ:~_[8��9Ϸe�D��wz�ܸ�m��tu?�T�[%�B�K��m�5����5�����;��>\���T�u���f���f���>F����I@�cJ�;�;4�m�Z:�Ԯ?�
ǨOz�3�esF8n��c���8���'�Ef���;�.�'�K�f ��D�Y����1���,*�Q40� o.�5ś���o������Cs`��.AH� ��v{�7 1X��Z�Sɻ��#���=�H�9�Ǚ���聂�=�j;Ԕ�x�R���C+���͟��w�K#,\#�&�**^��+�zO�׈���1��d6>���dڤ�F��������1�2UT�xc�8Sl�U{��K���f!ǻQ�+�����ǰ�b�X���'�W�SE�1B��I��86�^U�=����h��G�,�!Nh{�O%�����?zu+~�d,k�&ރ�b����f�(O�hz"��1��4�7z��.��~�YH�0s̆p�
*�ݸ��#���[)�)p���}7@�Bs��������V.;�����Q�`�Ha{��Lw�C�Qg���P�EM�<R�`��Q0߫i��@!���7�r�o���J������7���x+��4�-G�|�0�r�!|.
�{�i%؟���־?���[$�V�5�?/�yo�QrjX1֒�͎p���rk�kx&k)�!����H�qz�.L���΄���m��V	�vP�T�b�G�T�e�@�ċO�(NS�(���MP�,p,�@�g��ʟ�O�R�� ��L@�$-��R�B\Ҏv~����$�>!��*��|4���Fx�/ކ�Y�?�Ԇ徏C1~Cwn��.����W��jT}vܣJ�	 ��x�ޯ[{?�v��l�`wg��,�5�~LuNa�RH�o�	Sí��=%+Z+�8�/�uk8F�X�e:��t�a�*Q�S�q�xEtaw����[s�R'���@��52���:�{j�д�c���*N�gD +�6��+��5�vo�t}���i�2:V����f���@�B��c\�%o�oshuʡݚu���I9��vkI�9�y��x��<y8�[<Q���YiZR`Nb���O�`�S�$(��4�!:��o�	ҍ-N�,K�^GNM[��p�Y܍��FX�Z�i`��y��;�{6X��GG��CbK����T�X�$�����U4��#؞����B������.��⚞�MZ�L���X�y׎,��4D��_��hP-8��Ŏ�X�(|WǬ�7(��F��H$��*%v?�����]����'HMH�,O%�K�N$u���	�ƛ�8�}�������~N#�^�l�3��%#�C���RA�^��nز8������җxk�*=�P�d>H����e����%<�p��jl�p,�e1c��W�xe�6�K����e�ջ�f�}*0|L=`D>�����e#"��(< ��&����2d��o���k�\�R[��pl���V<A���Q��^�1�#j��<Nt��ŧKE7N�M�pR�
i�²���-��i�Ӈ��qQN8�-���>$�7j��jby�$�4v��#O	�f��\�v� W��>�a����W�&�����f5�~8l�R�����^#��� ��Хa��X��:��K�jɯ2���uUMC��
���[=���6X�֮�O�����K?3}����l ����̊�3b�[�"�ة�DJ>����}%
�Xl�|�Z�2��;�� F��߆�-��%��,�UA�i�=>�(�D�ȥ�I��F;N����7wN��P��L�hw�U5l�"�@E��%3Vr����ꆠ$�2�ttq�IL������c=�>��������n�7�����3�_b��c�-�V��V��	8����qmS��A�BeԦE����:7 �_q�b��O)��)���e&��rӗ�&�l8�;=��X$3����B��̫��`?�%s\�q\�8}�K,nWly	����g��P��1)�L9��X�1�64�_�,hw�&E*HW�;J���}�?��92g͎�;�.�肞����%àڀ8c�b|�E�`�.bSO �ce2����%��ӫ�7h�O+��-���Nа�H�N�+ǰ+��k��/�o3k:Q���m�3C�ŧ�L�Ri�E��)�$`l�A8c}xч��Λ5�l��Hj�w�?1%�F>P���X��B<������?y������$���W8��+���!J����w��ݸ�}��.�tW3;�L�^i�ԍKf��j�j��e�A��j�XB��˲�~E�Fpn�pis]�L=]�@T;����u��-������xiE���gؗj����#����A��W�s��U�f#WyY�������"�V���X7�S��Ԫwo�r�u�|���f�3F��d�@�M!�m�N�>y�$��lTh8�_[Hö��/���0����([����/�'	�z����9����udŻ��������i�(���e? ��)ĉm�� �3� j���{�J�T�yOӳ�a�����
C)�3-t˃H���ˬ��v$f7�Vk�Bk:��HK�vL
.��1O0�"��UgD4,q��ȃ��@�~�� ����k�9nX6��&�l���q�T/��p�\�ӌ�z�/]d�f�;q��-�v��{>��$7jZ�kw������ۣ���b���VPF��Z�n�#d�������@RS�|�ɼk�
^�;�N�LD��R_��d��e+dۥ��j\�0�V4~�6QmĻ���h	trg�3u��j�	^-8�
���iFkhWMxT)�������7�'�f,��[3PSۿ8�G>K��~ZT��Zr�d�?"&9h��?��h�.һ��:tfe�9��/�PU��RQ�߭r�T쟸
�5��w�R�]���RY��Xe=�U:Z��IT�o��.K@Y��bH\�' :GX����)g9��̭���&S��kD�;��RE*��2���~�����2Q|��U�$D���`qփ-��gM�|Ҧ�z4S� �YzQ�:S��77 ���Ƈ�A��Y�t�݉����f7N�'�O ��F=�����ݜ|�s��"T��զ%�M�b����_�o����'bK��,������)��}X�>��2F&z���m�~���IJ`���CkM�n��.�9D`�+(������P,�R��7��#�9�{B��\S!��=������W;�RE��"D���J@wW6wJ�^̪��D�)�.W��!0� �h����M�.��&���ࢣL�D�XH�,LͺV�}����?h鞕�7�r6�Y�f	�Վ���\A^�1n4T)��S]� ����������)���3�9r��-I�;��֑�D����$Z3��2��yo�
�L�����N�9|�*��Y��B����	px##��5B��˦��b����Qzy@y蕢�楎��u�B����ՠ�g�m�IQ��T+l�%�)
�L�~�`ӛ�O�P�$�I����h �#e�i9�b'�����MS����a֑�����$;��u��6jM���vUrDם�2\��ږM�|����`{\�g^�A�Z{�/�1k���2��Ŵ�sN7��ڇ��4�����-�.<��CH��ħ��Eg�R��f�Cb'�4�A�5>Khhh��(���P�Wo��<����l%��JR�~eڕ/���"��b�����&�����O�D,$n�yם&.�23φɐ�G�*I�L�P�3�u�P/��,@�?��u~�_���<�#�k��O2��$�k��f����ܩi���6��n)�]�AZ��3<��0]�6TX��b� �㎩�������褧��<��wz���QX��W��
$��u�������%��s��)�g����*WsV\Sr�x�1!�����0]*��$�p�E���)�m�����9DH��s$&<�;����+ 7�����ǜx��>kτf�>XB��]�hx@�LW��'w*�&��U^��i%4�b��]e݈����&#�x.��cN5K�I��=H؇�l���q5,������H�uY}K{6�
�p+�F$iH����ﾴV�WJ�>�g���FQpafs�p4��$W."'C�tT��TB�lۣ����e���T�:���ݶM���D:^�����R�� �q�[�G����ܱ�eC�dh���g����%����-�3{����P�k�Q^7����4�S�	k��p����t�{Mll~�hQ����(O���C>�G��1D�R!'���Z���݃����t�Zn��F���03�����G����-�[����VL^Y�� ���z��Wb�ۍm1�ߜ�� �=0�R-m�$��y��Gj�"~�͵�&�[�<�]�V]#ږӓ�r�va���m=���xl�u�]Ԕ?eT�`mf�"q�>O�5�q��.c��O�
XX�t�,�=-����.GC?�ND��X-�,�%gZ�A��θ�o�d�izi�ء�A��� �W�,��H���WE�?�*'CqV�t�@Lr�>�	±NH���8��ԫ7!o��@�>O�����i����A,�	�m�K5iV��A79�6�9>����n���~�īVy;�hC��I7 �9x����o5��������:���5�*�N��Rc)�E:#��Ta��A�4��e���3��RxZ����z������	��T�
9��I/`Ѹ2��N$��p�<R��W�@���N5�OuP���MC2KO��};	N�1�hx4Ϙ`R��c���u��O�a�cAz�T]Y_$x!G>g����Z���\��k^�4>��ʐ���E6F�Tm">DNGe,hK�z<�h�Y�FӨ��GW���X!��.��Z��˜��@x��,ƼՄ��[�yA���k�
x�*�],Hj�������6e�C�֛�H���yKP�*gE�t<��s�b��d�]�7Z�O��m;�p`T8x���M|��6�udu0��,�51��(�g�o�W���~�c�wx+�0-��� �?��a��!D�",������[H˞��p�zk���B��f�V��@X�ˏ ����������+���|�J)�?��� 9������� gIV��3ĳ� @�_=���?z�cP���V����ܳ3��U����x(R��%8��=�\�?�6�b{D-�`Z��(��}�a�e���Gb�8RFj����4���HX�.,G{�/��
����<*�g�6fIy�h��ݯ:l+�3��?~��:x�Y�-%�e�o�ޭ��P���c!��
^UA3��-W�#-������^��ϦI�~���Oa�m�	$�1-ݤa� ����9��Ӻ�X��U��j07�������皵�` �j�)�ņ���H��<�o	pLX�^���I<�	���;'rT|��9k5��.�jɢ����g��g)i��^��<�{4,u^ˠ�)_�*
!%�`�t�<ie^�}� ��Ӽs6�{����&~d�
G�oH� >"�-duzF�$H�_0@�'}db�_?7�Rq��T��x��J���k��'�nr��ʈ)����@�r��n"�|��J�F��%�}&r(Ւ1)�+A��K�$�r.�X�%Y�F֫h���|�2Nߣb�1L2d\�A���\���#�}�H��ß�K��X��IeB]q�a׍<��(���9�S��0d�4]�N��3�v��ײz�#Q����poTrCo�'��;J���lq�|����*���6:iMPA��M�E�c;������N���P��[WBX|�*{ךҺ�S�g�2�~��6#��+�Zc	�P����p8�w	4=/D�e���8y�:��4&�#� �N� �h�=����)����`��S��d!��|*�f�|�t��o���n�  u�K0F���O��4˽���^���8bxXpU$�x�����*��A��y�Ja����K@��UP���8}q��y	p�$Z-SK��O����)�!��!Dk���J�#�ě=���V@���b�]�#a�8�Qk����0L^i�.6��5N�|�"�2���>M�#���}�Ht1�;&E��xl�ge�$�2�)�66�����Z�^͜	E��M;E��)EN�'5�g��0�1/=�[=����}�x�G3Ҙ�i�9�?8V	�� �X�R�he�s�]Q%��sˑ��]yssiT�bR:f�C.�sRg���J���m�,�g�vK��	U�V4	��\$$�YW����[w����e=� H�cօ��������5Z�X&�����D-��봗��M�m4��s{d���RZp�P�"��:�x�DMA1����΂����* � -��F��,q��������p=L���y;���6�=��
0�Β�ЍD�������=�
Fe�_߉幈j^8�-!w�?��}�����+�����G��p¢z����*Q/�'�6� V�(b+�qω�BBZ�f>�j4��6%IEi��F�GZ).v����X�ÜXO{{��'���-5mzSpAVLB��8b8�a
��7ó#v�Y��!ә�rrV4��β��yk)���z����7��!(��� C��̼p���	�uP����S��;滷��PV��/��\k���*�R��c���g�}��s�9��Ѣ��~Hǹ��Y++pf`{���}��i��'�{�K3�����ؑf�.���a l�g*K3��DL�P�1
]�+�H���(��V_4�ֳ.QA�u��3�K���$4���<�H�8�zb�����Z��6ٝ�����:t�kW󦜏
S��F���@�@�w�'�T]��X�Pd�&�ǆP�N����EQ���33��v�RY�Y�]_&ޡIipݸm���b���t����P�{맫�%����{ꗩ�q���:��C�0��8Ƃ�c�i��Q��z�C3&�қ�Rj���;%Cj�!=����B��n��g��씴[��l�mV2=mfNH�#	�/�ɾg�E�E�+�<����EW�0�e�ʬA���ˡ�C������0����o�t�_H��*N���;گ�=��N��J<���:�0N7���_��l���y���$����͐#�f�_P�H7+8`Y9�v�b��:���c�:��j���l�CEc&0�D?x$��`>&M�MտN��9<�g�2X�|p��}����TʼlZ�9�۴�as� @(�ǘ�	��/�g�-g�u0g�sŀ4OG��i��p.01A�:�����Iqd�����s�@��4_�"W�Q��9�5�Ӡ���t����K�?�
�����/!�_ӊ��Z�Ki�IY\F ������Z�*�[�Yd#����i5�T�]���(����sǮ�&V�0O3�g��1�2�R���m^�
5��>���wM-~�_u�<��q��bn#��D�]l6 H5��]t�AQsfp���;�L6�ͺ#�\�6��#�r�Ɗ Z��O����Ny3L��H�]��;�p�h�FG2\��,�o�2j뵭�W��֯LQ�a�`,QٱL�ɮb��˦����.�����ד�~�	�Y����)8���h�Jpz�+������*J��_2��!C�Ϥ�r��9-�j���Y=��GJ��)�ՙ����F��_O�Q���= �����_���L.���w)ME[���~R��V\ϰ�h��@�a�5&��!��*�i��6�����!��ۥ}�+������!�y���G4�{��n��qX�qW,;�����2tΜ�����*�ѩ���~f�*�:��?�J\Y�@ֆL 1S`�?%��,��18f繕~��L)]��"��b���@(�l%��8�A�8[FEs;�'����6���nuB��1f�����LE��vЇu=�s0�;�炠��³�
���5o}��"4����T2���^��e%XV�-]�|�I�W_��!u����i����1�x�ө�Zi5��[F�����_���{A�`;�M����f��Vxn{l��Riܚ���%�{�^�&��i�ZY)J��ۧ��
���s�������İDt�o��X�����-2	�>z.� �ze��'1l��
m���Kk����~�ҽ:�E����V���te�TALX� �Y>Z�A!�\5�hr2�KtL�*מt���Q�'�sO4��Hl���v�b�䴚���8�f��L�
.5gW���-ӗt�w�����Q	k�M�cvR(ًMu �fI��h� ~�h�9�`�u��L��%�d��ц�e��KP^�~^Xr27����?E�z�������0�J���.��S+�����wR���p��F�]��܏e�:�D2�	�)����c�S���
����������m"�'���V2�Dr��8���m:SVkX~��S�A,L�"V�c�*��.�>� ��Ds!3;��8����Q<0k=�b��z1�	+3��֔�HUȐ�U&��m��g<>7���JC��-�`T�x%�V7�;�
3/��e�����l-(�����A<��tu�JU>.vjR�8
�|Z6)d�y�������cp�
[��c�7S}�\Q�w���g����梖1d�>����"�7f�.���T��Ƌ�5U�²W�MD©*��V0���m�ͩ=��f��k��$M�W���
��1����6��*%+�T��ﳏ��O�K&&hӀ���5߁>j6IA�Ƈ�~۴ŵา�>4Sd<���{��k����t��dw��M�s��R��lX9�G�c��A���.�$-�����5��Vᑡ>�(×������Cu��NR�����'}-���h�8kM-�֝�v>�F/�Ɓ��K=��/g�9_0��ϖ	X��,�}�̧�̞�E����,d>�Ga��1B�.#�T�nX�.B\���>�lu��SfS�T�������1�3�� �mZ�F��s8]�Ґt�m��Ns��*���22�p���ҙt�!
ki�����-s:S�_#Y���WEogZ��;�8`}��&D�q!BS|��Z�Y?�-e]���P���K��.��1Q���wQ:Y�[���^P���
�1c��`��t�_eЇ�S٫&m0���^G8P�E�<��4C��,ܬ��)��qX-���J�^�HjQ��ǉ9� �._����z���BR>5L����l�N��l��'���Kx�(g2�_�ˏ^�������2j/�Z��n�D\z���װ�{�؞� ��>�#���2gE���m����LBL��Lf��g��.�҂�Tcݔ�z��V��,E��W���E�Sb�����vqA'L-�b\�̮���4? ����.3&�Oe��M�7K�����S%�=��RU.H|>I���z��Nj�&�?�À[l�����Ĺ;��&!�ڣY��Q`�ϐ�T3�Y�,I��@��g�ç�L;HG��9iV�E�⻹�6Q�J�N�d��R��W����=]8�3(4$�EQ��x����D��7�q��d�E�/��E��J���S�����h�ӊ�wP��2~�N�;n���>fkP-�KS���dEH�1c���1q����n���A����f-�����$���O��po�H���h2�o��:s �v`*�,�u,����8����c�_�[?��+8~�+]��!��W�-��B���.8HG�G����B�͆=���B��͚Y(�>��m&�[�%h"<~�w1u1��a2��4ǘ�Ǫ���ӂ�j^+��{[dU�g�JHͥA�0�R�|N�]�<�8e�\ԗ��"�}��[h@lĢ���v~!<�X��m���
�1R���,H��,y�޳j���׺�\e��<���%���*PK:�|�0�y�c��MGT��X�t�5�D�����Vwd�N�̝�_�r I����xk�bƑW]��f���U=r�}Y<]<	�o��Sb��� *����>:G�|]����;.~�+�w���M�#�����~$7�]�e���)K����@�*�Lf�=_�z���:B$����4�^Ǉ�cir��P�GֈM����Aԡ�ۚ�����]��f^N�Й�����D�|L9�dKۏ_4; >��ĦJ��,��r/�<�	4�[���j���;����yZ�<�n`s���<>o�����ci�wjK������K�w�[
�1�G@1������Y�����Ƕ�F��ԩ�7i�g����(��le��9�l%������฿��,�w�:@\��������1O"6
�������<͸i-u�RC�;�TA�X���,��|�ke ?ڝ��Wu��1�+K�r�tV��8���51f6�u̒�M��~f�Rp���^��[w_M�@�~�����R
�L�&^���2�kH�ǭ�$��;' �^h�"_(/H?�ašӓ�!����G8FM�n����cM�~�n�=��=(��C�~{4y#������ $�!%���o{�I�7)uC�ѩ\B��k}�Y��HQ���
3�nXGu��<��� �^(<�Chd�k�#��2�����W������y�����5�r�_��ֿ��ў
����Ơr+��������"T&|�<M���ʃ����q��|��G�O���X �X���0�E���5[%o�փ�2+�Ȟ�-=�����(���g��ڗ1����u��?�=�c����`Ѐ�E�N���O5��B� ����Vٳ���I��u{*m��β {Au4��I'֜��=����[_]vos��UI A���fA��@lc���t$�@9l�yW�y��z�����Ց�����2ܞ(��L%|Y�.e͐#j�B��i� !ʱ�$���^�lmx�D�9�IO�Kh����L��/�M{��)��]��y��t@#W���&�9����Ȉ`�Kg���Ğ��S�KbD� ?Q��(d���[k�_>�E�Q��pba�ݲ䶉����Z���/����U8,sT�����nY5Q�O�RS?^�5��ġ�O�槌�a����%, �4:$:�O�a}7�K<q��{����.T?U�ӗ���_��ty������F��#��<�Z�����.P�&�Z�#@� �y�e}߀�9���.��EZT�J[?8R�"p�o�W�b���؀�DG�=�8�fh�����ի������1m���/vQ�֍�<z��T;�9��~S*�+A��I�y�i�c�"N�1APC�v�B�)�����%鿸�,�k��(j�3{��EȳP���	�R�MV�9G�M�CUd�Tq�tX�IޟԠ<h����V��*�">�9�^=��y<��,S1'�l|��1���ޤn���fA���'�ω��ѻ}�l�#,�``��T���ԁZ�?�]�BT����D��jK��2#|�4�B ���!�T� w��Q�~JN�X���4���k��+�^�	� ���P����[����v��U�8�M��w&�����@��a��5�7q�G",WL�A�sXmNi�|w����8�%�ɯ�p�`�Q�j���t$�ϩ!He� tm�G<�I~L�r��>�����B�)�M�+4�,럝>����&<��to.}W��������zb�`�+	���vy+�n�'�4�]�1\����N��6�M1-��82JX�n -�3��Q��נ�s2���?��UF��p������e�v�2#-$6�|���[�.���%�`P�A�ݦ��i`���%�`�O�(�{��g���� ��t�h&�s���n��&
�&�+]����1��l}6`��aGS�S'!oe	��&A9��M�%�d����q���iN\أ�5���7Cy�D�fO��$���(��sk�t��D���׳�t���G����z��i��!�6#���7����գ�/r6HOn�v䑗��LT������SN`p��5�@���ҋ�݆�}$�l�!��Qs%����{���x�ʱtyS�먫яq�Д����rG�L�@7�W���]@�4J�^Ь�]�FT`�T�Ϗ�U57������$_eC�Z���� /"�+�ѹ))����7Б��tYf�&sc�9��%=�Y�[�\�	 'Y3%<
���j��C��߈M�F���e �V�Q�����s;F
��K4aRTQr�~Ni��S���Y�G� ~�Y��O�G	�_�t��XޝchݡCx
b�ch��w�"-���5�Ŵ�.�Wm������v��d�Q�%y�щ�e��. ��)�ӯR����=@�p�1��=S:_�[�t���E�#��w6��23��nL|H|��W�S�#��f�ҳ�u�ri�jO�z��}��-�گT޸�=�&�Я���,ٿ��	�[��L�c�Õʔ�RlU�"��.�lP�t0J��[o�Ѳ�mt��#>6��/Qp�5�D{����<M�W�pU�"R�q(bX;|.�c��@5�{�ShV(�H)ߋ��l�ܨǅ�%��uY0��@j��#W������xm����a`y�fx�ުDyދ�,� �q8�L56)��:]��z�Jqؽ�ȍm��ah��S�)]A{|;����o���m̃�IS�%�Y�����x��w��Q˷���&!~�g������=��J�|"#�1��ˉ�Q���ɫ'Լ^�����1
M����4Vͺ��	-��ӊa�:��$�X�����2B�ACQG����Cn_�_��75i�N] ;���1O���=��en	����"��6$hg�����������R��9]�d�IuЈ��:_��W�4��xM���d~v:��u�-��ܻ�2	{��K1��x� ��m}XӮ��xd���	ع��Öb�`p�x�(j���`���,��z�f�]e��}2#x?�
�(U>�5��u�̬�9y��Eۡ��T���)�|Q=��Kٰ	;Va0�G��f�rA������aj0��: ֜5W�}�X��?}�]���f�B��%Uwc�:C��dE�����D�����N�ut��=�ƺ�����8��id���񋄗��ª����9s��g��
+�[��dA���M�v���Fn��7�V����S[j�H��Ö��z��������n�(�W�$R�$10�o�����op�f�n�},��t1�x��:��x�o�*�b8�\��&@���Ǭ�@u�~�+��T�Q�V�7�#��u/��#_#<N�����Π��u��.S�e������J����\�P��X��x/m�/�VG�Y����%��U�ơ���Z����� 'ߎ"�4�W��-.j����E�������,i�q���,[���5���*i��ݛ]��:]�A�aQ���4BbS�����	����������`��%c#pR��S�O���1 � �!$�gLc�Ô�j[GNk�]A0j)uÖ�g�Ю[��[ǥz���S"6R�_{���U�T'�׷���kғvM'0���?����{-Z^acb9Ӕ�v�� =i�̵��Hzv>��pY� ��f�I��!Z�\�~��D��|�9I!����ڳ�a6Ǡ��WFΈ�b�d��B�Ω�l�S�Tj�e��#����hӒ�B:j(��$b �J��a�>ZH]�y�p�5��^ X{��84@��l%�ٯ�W�G�����M�)0+쒢�B�qt*:��c�
��W@C�K/�"��'��If@lb3��9[̂��=}x�����o�e6	�ok�{��q\�p��ψQ���V�8�U8Cҗ���C���z'S��NY��(�1���Úw����3nK���ƴ�֍�B%G�g�N%Y
�C���JA�7��ʢ��b���f.�%��Uf���ٌ���b�?vٮT�L�&[�+�m쨸_�����KܼxHӗ�ܧZ������F0�n"+P;��(�Y���S��Wyr8���y#�T�`��q��5{��o�&�直ՙ���d��[a,*�;�BFB�m^bK���!^{$W����W���*������jmr��<�s����"K'
�J?���^��yZ!J���{��@Dz�d��x�I���S����9<	�E�jޟ	��ӧ��NN�A��F����|�E;:>�+#�����!Q����	ȵ��|C�
����-�uQ c����{����c�+��r��6��B����|Eڣ���d3��U�J�]�u�ӻ�-L��W��u9��}��(�����j7[-��w@����V�ߵ�b��=�a�*����tx�U�P랓۸��`�@�K�ksJ�3[�r� ��ۥ�>�=�*H�l{� xB�"#�k��� W�V�m�U�C{�p�7Q����6A�oˇ{=��S�1���$���?����7��:#�8]���7�|N�g�������Er�	�����d����Y�T�B�c4�i��T���ڳqVp,����bφ("U��>��mRj,bxv�:��c���"="C��q��;/�i�)mH ��2�nS{j`*��}�V�jVГgMK�1��[�8C���x�SW+6���$� ��ءG}�k~�j�� �	�4�Q�
�����=q5�7��#��-׿!���s�8p�y�b&�64&�Hc������-�9D9���n[�	ˉf��i����nxBY��ď���(dWi�u��LN(\ye~�T��mkӸH�I�:�޼�����V�*}+.�}%�U:�����nϔgװ��?�a��ݚ n~�`tC��˽A^�8�,4e�{�Ze.���C��*5_��q���u߾m���MEYZ^*q	+����Ǔ2GP���6(�m���|���Vd���ҭ �m�wlΌ�N�� M_����C�����?)��W	�1Pա�`q��<�l"g�����!�s�@�[�5�υ-[|�I�q��[�y<�z���Ho��*� =��e�ݩ��y%oI�T�#<
H�wY�_\�ן�gO`�~���o8(Z[������Ӌp��m�G-���i�{`&���K~���6�N(Ps�7e+�Z^F<�g ?@�������(L�o1Iw�}�w�b���YC��f{��כ �6����3��"*ԡ^�({?x̦fW�����9�cH�,��V-G�?���$�9R9��A��u��n�;�br�U.�HW���@/�9�JT��[�Ͱ���B�l8�ܾ�!����b/qv��,��^L	!QG�=�/�� ����zV�媡�_g�o`}����������/�=h�;�[c��X�`Ǵ�|Tn�d�}�x�~(R�W��SaT���~���A�@3	�ļFy� 8�����7[S=��g��tKo�|�� ����+�Lz�%[H�K���7E�˴u+�6�������͉x�wGW+���I�Eŉ�@"hxz�2��(����p�7*%��B�W�����VֶNɛ��N�$b���C��U@�t�%�d����K�+.�Ryq�7�iK�8��%���G�H����`͒W:��?�{��
9A�+/�M�ݿ��:�9Z�����h�f!V���6�Ӛ��*�]�/;(�S�w��I'A���Z���N83�Ǩ�{�C�����t
��E��2!t6�l&Ǟ�մ������Q��!N@Q�}�oI�Mf��|���O��_�1�h�#Zӕ�[,V�>X1����cy��	���("Ӑ_j�v
A��I��uU�-�(��Zy)�Y�����������.z�-�A��ZM9?̣�^���B��j�L��L�i�4
Yb�V���(n-���R��t�A?�P���)Զ�}o��H��6�}�{�gO-�H҈�<ɠ�Ĕe� �\�y�]R4�SM4`��A�;X35&�|S�z�_���H=�Q� �n��@8&�_�j
W��q��5w���/-R�j���J(�B_�̟��tM2��vu�0�8�%"=7��)������5�V�JQV��l��Ϥ-.�k��O� �J:�R�����	��0�I����~��Q%����d3!) ]�%� e���;�Ń�A`X��#[`�	�Rsa�P��YS�S��Q5�U�e5��\z�G�j�@���b#P�}F��K�t_֟���X�ca1]���8�#=c�U8Ŧ�@�#�6���iT��ʥ��z W�,�+��
�8��5���7⥭
u��׼R��-HU�F+��,~;�x�UJR%��s1�P�DC~�B�,6���-����&��K
b�;�Z���^���{U�B!G>9%e�σSz�P��gq5������oz��j���=�+��Xi�3F�˓�h'6:��vˢx�:�o��#>��r���6����M���������%�]Д���Ѿ^����![�1N�g��vg��
Ս2S_.e�.�#"*�p4�3&%�޵����i�I����|� r@P�K+��Mϭ5pe,75��'l��~(3g`V�RH�Ҕi?"d����}SdV�x9����'D_�{�Oѓ�6I:�Tcc^=o�ݽ)l���pK�d�����qz�,��Gph_\���HJyk-���ɤ�+r���P�(�:�Z?jw�,-�U�_��kM�ִ�R�7\$#&C�zYl�g�`zи�9?�f�Q	{|�KL�2*�U�\RB[�.�9���C�Y�i�\,e�+�s�t�!m�DRH0�dn�@�ͦٸ��W��2��E>[��S�m���%c�$\}��q�#�%�!uz_r(���Ȼ� ֠�� �����q}����G�j؊�$&��w.�`�&���e������O�sE�M0>(�yS�;�G˸��SD�0��GG�t�ͯ���7j�Q!XMlW_�m��B�D��:f4k��̭��H.`��!J.��_Z�)�9S�ݢ���7s/R�hϾ���b�����p�.�:@�X�i��+�3Y�Z�7Eժ����d�'�
{q���Q����be��=:vZ�ȑ��#�`}�6�� ��f�n�D�Z���%�)|4�ә� �YR���2�,�n��d�k4Q�.�'+��h��h L;p_%u�?�����6kN�(�)�#ք�T���i)\,�"X���v |�� ��]&�+3��p���� �Ό5/�B}�m8m*�}@��g��)���4:UH�w`�Xo@40J��n:��6�o�/i�J%�)t�f�?ASn�Ъ�
j-��^����>����o�����W�`9k�:5lB����9ۦ ���^�{����������G���@���.9�,"�pd�TR�=����-��g7���pCm�	m�����FS^���p�q�>��T�E8������B%��L&�=�\$?0n�ء��FQ�����z��] ERC�Q�5ldO
��:��M��K:�φ✙fف���(�s�����6�h5���Z�Nr���1 ��J���k�Q�g�vr�ܶ��@'�U�O�|�c<��Ѩ�TSb�X	%�;�'�F��=�Ä�~��B�w6�n��3Ԃ`��3��'��=�y�0K �)�jki�$�7� �q����CL<� �0��g������6�~��.��|���o�GWf�;�	��"N�T����ً*[��k_n� �Y9�^�s�f��E���5�@�W���ܮ�ŗ�-������7`D��`b)�Y�O|�٢��������{�j�L���P
��
k<���=䬩�CÀwy���Q�e~��%�k���3v^@�^-k.�e������+��dPd��5��9��4�p�Xq�޽54�F��@r�L���X�W`����rT�+�ق	A8��%WQ�8�H���O�!�ȴ�����`��;�c?�u���`��P��+?�Q��O�I]J��Z���4�~��Y�ü� �yC4{���n�������q�Y��&��yv��,WvP������^��B(��Au��`L�bV�3���	�� ��:!�[�w�UVǅ�e���?�������~2��ѯ�byl���b�r�=���  �򢵫�������H�⣮�.��� �/�IZ!S�}TD��+h*��}R�.C�أ�����3�(nb��:�����p>I%3���͚e��ϭr =���2m_AQm�)�Z�����߲��sѢ͇�vՕ�ٔ8���A�t_�[�!V�Fl��8��A_$qw���ybN��=-�]n��7�'�L��a䂭����K�����&�ߐC�AM%��yigWg�8��˲ÔMԧ���������"t��T��B��%��Z���:\�&W���f�߈�)͐:A���f��b�>S����QS�F0�����W��5|A��L�Ƿ1�Sok�BBT�Dj: Kg�˵ʃ��R����ݚ�@o�B�Nd��ΏbBꉆg2F93S �Z1tL\tq�����&�}�W؟Z���@�6�s�L6��3��=?��w�x�3]�O�
�3N��zm���;����E��V���m���<�y�a�Td]�%����d׸� Oe*�#�	F2�k����&��'[i��cRGfRjV
�3[f)w�EȄ���졃SU~�$�(DX]O�Q���j���\J��"�
<Q ^,�q嫛R�x;к0��<�T��#�W"�H��OW-s�#8��e�s���8~���|n���P?��a7]��Ck&d�gOi��(6p�{�a\]	��9�n�M9�y��͑�L�A�߲rn��+W��HB��
�Lk��+���$��'��\զ��ƫ�j���X��Y+����䄢�	��D��Ҏy@�K���:M� 4A��d$7�55�Uý����2���MY��g֚r�_=�́�th�Q6�O�UXZ�V�����9Z�@����x���`/���V�{t�qXd�|�+�&�1���(G��P�L�>2+�u��锭Qd���N�:J,�[5����@�3�T&�ݶ�w%5�n����E���u�V�����6=�1e)����ՈV��ȼ�a�N�A]a�{�C���7g� �VeZ*b�S�b�!��ܫ�Um��R���G*j��{P��sĪc*1�g���Zǁ�ZXg��bi�la �U���r���^x-C�<Q��z��y�_�%z���+y�k����b7�w���x�fn�x\���^Vy�{�_�R"i��P_��`>���Wg���,��S%B��Gxcy��A��-f�uu�V�y�t<��WT�p�*R(7��fj�ָ~�WdZ�mH����Zt�!X��?�����񗪹2��
���Qv �l��Ŝ�JU":oܩ5~\,NatA�K�Ba�>���SrͻTS�_x|��Ѝ���Ya��Zep�b	h�{��� ����=�e;��S�G���9D~d}��XIs� ��`?�z��)��W���T^(?���;��-BE�*_70��R����ܱ�ҁ�q�@�3�<�C��VTS67�����;Fjl��ڦ�b�J\b�}��}"�h��Ŗ�;$&�i�6��?�u<~j�������QȈ�K/zv����t��zY�z��s�a6���g,m�置E�:S~"ž|>��vy��njbd x��R��6~M���Џ?�*��U����C�o�i�|&nh����7��xk�I�.��>��W���ϕ��0�7�����=[� Z�_�Wn��
�Kg���3���F�w�����w�tȶO�"�%=�[n�����-��V"@�/U�{���Ob�sZ�0>��d!�0�ω&� yjQ��h7�|�{x�0Cai���c�x]������|��!ρ�*��Gb��ߍ �m�76_��cs�s�+ւ�̪�\��-e�Q�֌.�t֍���u5�׎�ҟJ��4�;���S��3��'ܥ�DVps��,3�<3�T�j`Tb���n�ߖ��d�P�\^�?r��+�	���C/�!h�@Mx�XPt}V����kP��
���u=��*�ڇ뀃���&TFuXvZ�j� �����D�ʸ3����eg�Jz�c�)����3����J���c�����F��Y�r4���S��e�8kh���.�j�#��R�:����� b˓@>]���b����g�I�e:1j�*|���. j��+e��%NZ���~�a�`^_k���#[t�+p/�~`�]������,-p��M�o�O�n�&5��i!����$���w��"����ơ��-�F���B���#OM��}�L�W�PE;�m��jbr9��Qs��3�_�Io�m|:0l:�5u{T)|��ٮ6ș�l..��I���ޣ��6MZ����C����R[����$��`��Y���&�D�N�aۼ��k"]��b�-T�|��: �8cu��*5q� ���V�^�aRg�]�w��j�ZT��|@}��D����k>��ц�d�����I�^�!
���BylJ6���'�~��Չz�\��Y����O�Tۅd{x�����$�9�C9���>�
~���A�┭f��_AmJ)5�s�뢀m��v�ֱ�#P8��f/A��d ���rn�J���T���?�٤��$HVV��q��j�F�Į
��"2'�3��Ժ����Dc§>�{��|�� 9�Ѫ���B!�Q.�P���σK������P+���w1_�z"Ʒ؊��Q�:F���Ng8��
��;���7�l��|?��Q��5��@�c`�) |ک��|�TD�-�ũ��;�Ln����z��ܮ5����'���`!$�dLc[���5��Z�L�94w�-�d�iV��d�j��N�M<�~.ӥ�[\x�8&�c�H(e"��v�Q5����ɪ/��0�]��j:GHܒ�o�L� �pٍ�3�>^N�X��� �q�ǴeN>؀}��X쪇,��*�;�m@�	n���ه�8o+�V��u�y;ok���7IB�?����jR�M��_Y~Ɓ�����'����5z�01�^t}�Ҏ�4����}��ZZ�}�f���C�cZ��.[�Yߘ����\�+[Xf�K�$&W�I�^K�[[��m��{� ��8q)�VF��zH��<qpjq�b͂7��j��r�U#�ֈ� c�{ȷ49�f��ٿ#R�uWU�����^�x��D�e���0�}>�q�*�+ Bc�M���>.(o6�/D�,pP�da���,�7b����\!$�X`��7�@a��D�#M�B�H��g�i?H�N��SR���[5�tii)�R����L�iv�${-������O]�y��B��V�S#}��z�S�"2�7�+�^U�{f�W@�����|��5lōR�߬�f)��������z��he����ms��/��Y�A�d�G�ͩ|�i�T�m��Y�#�d�|��e�@�"n��nD�y��&S2��,M.�џ��+H1s�хm��	0'�?�5a�<�9��Y��1�I�G!�V0�)��IY90�Bڠ���%�'<�
���l?{�f��%E?�T���#�8Y����� �^���3/On)L�S�->�#*���aTP�#Mx&�960�7��]K/����D�ۂ��@\qJ��Z��ˌ����n^�0��\�bpM���u�����"�ܨ��s�*�r�1V�L���2��h�	J{�\�3�S��{q�1���}�O_������
�E�nƑ=���K䍡!�+�:�r>A��-P7��X�U�!Ji��;� �swƧ���=�Y�`�#4Tw*@�kx�f�Q Y(����8%��9+�YYL�i��1��z � ّ#�g5O�/����Qn7��`;b��l����E
j��|�mcy��5��F>�_���BCfUsdn6S��r��F4 R�e!��[8�)�^nrVK�����ᑊ�]�k\�c�P73�[�xO_�"N�ʺ��N�ZaK��ݞ`��n���JѦ�C������Y`����}�[$��HY��n�t�U�u��j��|+'�N��ĲC�EV5 �h�c�+�/(��P"�$*�t�s�L(V8�(d a�w���N�"��2?U����� ��6�kY>��e��g�ceMCa5F�+p,������$R��Z�y�R��0
N�/���q3�޵�i7b�w��[W�G�|ȜG���F#���&�)*�ry�M*+bQȦ�''~U�d���Q�><��L@�Q�,!'�R8ȏ�G����_�
}C�q?�[��M���yR�^x�e�\��/�C�d>$Pb �hd46}�ѭ��� �C�t��_�!4j�c�Y����`>�Ge��6���3���'��$|}�i8��g�bG�+�I^���b�
rj��5{E�0��dM)�n&`�/�H܏4�;W�p'&�y�:��{[
���):I/�b��o��*&�x�(1�-_a��"d�S���`���_T��PwB=v��ώ[���qH��Jk���X�����[ً�wn��B������Ċ��~��x;/�-ӞL�Ӭkw߂����Ҩҗ7N�V��6��ZwNOeG�l�1Xw����T4E���#.�/1��V�B�IO���(��`�i�!��G�3���9�Iyq=]ɶd���I)p'&UP����6�m�f���+,絻E�_��ء,I�$2�W#��� iN�N�( �Qe���N�S��w
�w��9�kC�~����%c�kd��w�S��	4=-�	��a��Ѽ�N�ǃvF �� ���oP�Gg@���k��;3I@�(��j���X}˘����ͮE�;.���g���}�����ŀ�]��o��P�2�"��Jt�jl��]�𼴮���V�!H/�C٬����� |��0���X���{���?�%tRnd�$(�֎C~��������./`D���z닿��XJ*<���<�ǣ\��<�X��IK�Xʧ��w����Vwh���A���\��.'���7=?F�$񽼿�\<)b@�����?�+�`�,m��#k Ub�%�;&y����@rP���*�!H��_�(rz1V�_#!�i�a��j�?�F�3 C}G��~�?����ƕޏ��!S&9>w�fk�Fx�R��`������4-�h�����<����KXr�xn�f��a�d+��)e��V�!F�ʴ����x��V���a��֨&��VՃ��������.����<4�Թ��;G~�hs�h��y�߼�(��������յ���PQn\H!�Rm�f���:J���#�YZ�S���xap���ϋ��Ø���]$�7yv��p�3���/[��Q�G�C<��X��zg&Cn�i��K��4J�6_H�j���b`��V�۪� t҉S�����(˂��}���6K�&O<�]U;q�M�-�� s�$�#����(�az�cܮٴƿ��k�q�+ӫ�yI}Ra��w��O�<��//Z�R�9�eF$"�� Z{+Z�͸=�����1<�������j=h{J��R���޸i�DJڑ��_��{�!���{P�R�rZ��K��R����SJ	��MQ��~�p�*�1�vv�N��3eV�I�|R��M���qC��F��� �,o��9�x����B�@N��5��Yq��P~����K"���S�ӽO��J�p��D��cܣ�U�n��[֞$�����������J+�5�3�I,c(�aoV�*����"-=��b�I#<LB"1&uA��M��jp�E�8�h{b;d�~�|�� �
��;-	���F�B�aؐ�xwZ����X��P�����e@�N�9\�p�qX0�b�s]�W;F�!)<1LyH2э�ը��β��n���N.���gT#��YP���
�:O�9|�a B�upo=!���lNW��C_�Ht��-��y�a[[��QAQ{�Z�|�o��Xx]fp����Qj�i������y�)�s� ƻ���[ݽ��7$��n�v�yၼ_�9W���@��#y���>�����TM^L���;�t������"�-+@��@.m�6B�c��>˨��@� �7�O ����[D`a(� b�QjlT\�p����h��;��V<��pN� �'o\0�&(9������z-�_`�R�sr�ץ�7�7C�?<�[b�L2^�)e얞��u㸉���Q���W+4g�o	{���ָ3~ET�p�ӄ��L�+��U����S�4��(�����P��r�����pD �4З��Q�5��X�%�ot��H�j��ߋ��0��A�9�e`��E�j�$�V��?,�}C?�!@�W;eX~�=񀓀�y��_&���m����Rzz_Ǒ�Tuz���&~q�^(F�Y<a!�Fƫ�JN� ���H��h2W�#�����o�贽Un�CN��6����G��8a�X{�����y/r���ِ���t�d����%�	����Ҕ�G���&f �<�WhzF.}���R���'�Ҽ�t�%	��Ou�r���S�LA31���&�ƲwB���"T#Eysd��Mg⭟{�=�h5t����.��[tt�+�f�?�T�r|��̌ǯ�&Rڼ$�K	�7�8��=\�'�ޔ�#�\q& c�u�mN)�sA|#�߭vR٣'�#��# `�x]�˩�O]����p�~v1�8<@Q��yrt~SUK:�Z8SaP_��0ؕ���J���\�nV C��S���f����MK��w߆H.�f�������P6Do�'l|P� �v�o��&���`W6;};8�����g3��
���7L����8����P�'��B����#�m�Z��v�N�,I��۾�]np��T�ڰ�&/��v��L4�Wxg� ���p�2���=(W�(�c��bESK����85�:�-�n���	�h��P:i����� ���Q���RpAQ"����&��8e��ϡп/���'�^��kE���'����5��M2G r�Iq4O��^ I�ѐ��JW�Ф�� s���^S&�+��f���r�
�q�����o�@�p��������h�4-��a�pp�W��;i6��:D������ax8p���2�c�K�zg���fӒ6�Lz��o۬�i��Ɖ}���pD���h9��w����{���[�`���S8:����r�Q���0ȯ�_K���tl&6�ƀ��;Y}������YX���|Y悆B�^�99��Ȧ��\�q��� ���nmE	4�D��^�C�-���.V\��x�.
�k짇��}�x�RQ�.��7��w@i���1����8�#Ӟ�!M=,�.J}�H�h+NxvtЏ�%9�P�p�%O��j��9�9��JZ>`����Y_<����T�����~v���Ѫ1���^�	iYTOl��0�� ւ�E��	M�� 'P$��2^w<OCSL����Z>�I��6�r`z&B�_�	�`����K%LE7Px	���$n��|�`��J����j��Z	n���'�$�RE�Qˑ�?��>�
�b�W}s��?C�^��3�'Hk��Ll{�����$�0�&� }p����d(��9�RF�7iI�A��/#v�7�̬�B>W�&%�xTj��g�%x��D�O���G�,|���D�zߢ�$�t?��}��\5�YZ��qB�'�/w��J���W�A.������`l4c�@� �p����ק�����*PY����1�V�,_����U������}L� :Y��k�/�@��5�Ν&���S?y��f�]��$��I��Pd����O'A9ɺ�{)q����3���jU��!�.Wn��0cSq���D���9�bK�[�JIGT�W���0)�w2�< 1Y����O��������`�i�?<�������?}P�|�;�ux���o�]�-�-~�V�Gι��9��`���ׁ�,�UP�;��-���ڦ;���J��l?����2Wb��ZU��`۰�]��O��
�ks�ޤ�*z�Bl���|Bݼ��-��ŽLI����c=��L�l��>q���`(hq��[t_��G�6��\LҢ�4ݽ�8�B�P(��>�bw�m���Ҙ�m�����m��B(l|ѕ�/}�3�iO1�l��x�JY&u-ߋ͍qC���z�=�r3�/�s�nO986��A&��$�aK]�ʡ�f)�����1�I��	^ in��[�v�N��ؾm<*74U���h��f��ʄ�wXD~���TQ�����_����m�*�W�MfО�2�oX5Hw���x��!kߢ�t���d>���{�� �f�Җz��)e���[KMT�2��w��v�yڀs���S(�nO�_Vԭ��h�m���IF�� k^��)1���<�ႅ�����Y��<[�v���M��Ƣ�Ԝ!�@�-�d��k[�4�u���:�X��,tjC]󔲉Y7��:�4"B��K��7Bk~:��3�)P*s�o�ݧ�;ݎ/&˻�qK���ZN�`�4��Y�ܺ��jH�����ŋ�zf\�g #ɎNT�~���Ra/�GȤL�fR9��符��9Vj,۹*_!���0h_ǝS�Њ��"�"u��ď�gՍ�$�e�|��ѳ{٪kEklc�g^�<�)vO���q��X��YNL�^;����:��O���K׹��q�ؖ���nZ�ǹ
��@s�����D��>#���kSr�W��um�� |!a�5�3�f5t�+�_K<��сyI�v��ܣ_�$��ǭ*{ltD���E<typ5��l�\�-�\�t{8\���O�[��ߺ�)=)x`:�p0 �pFP��t��X��ۀgv+PF_X��!2��۔R�kzLʙ+���x�7Im�(S`��%���?�Gb�Y,�k��Z'J��b��rZc}���G�N����Z4�U������@�l�L�"t��<`��ӬTO�,Vtw���֌+]ʁ~5����ioC7��v��V~�OF�](znM֭�.j6u�&jI]>.��O���Ӱ�w���/���Z~i�A�J��0O�%h}>X	j˺�15]���nûO+l]����4P<�nZ:p��K����k1��8GA��'e[���׶?���F�٩��H���mL�+�짔K��*a�*_�l���)�G�.��^f�����T{�w��_�G�CY�}U�<��v���5��섙���K�k`�=�#��+*;녧!���%���ꃵf䃣(-ٮ�v�@���,.+ ѻ�P�6��h�q�^�jQV�|�c�D��!{�*��`Pr�CC`Z��U�y�]��4cE��B�M���T'��K܈.�h�F���aƆ �$9� waFķZ��3���1��#�]�ضq)�4�-	0�a�$�F)5��lB "`
��*r�~�������%�W�)�̌As���c�'�-TE���ڦ�A�GV���z�X�k�E��r��d7Է�9*�u ��Ϋ/��W���3
�M.QedP�dd�8܀�1|<v�sv쳿B$DXGc�#��bG��[Q	��i�Fx7vUS?�4��ܦ�l�£#��I�zL7s�������Y܋�?*��3|O��Cj�C��Dy��uNniO<��~��L��Х�����ɂ�h��f�)G������
盠�#�j�/�o?��tK&\��9��)�I�sR���g��YG��y����b���ݑ����"�[��9}�1$[��X��F�n�M�2�1����b+��Lw�w�31�^�T�V����{ox��kv�}h*|E��$���+T�՝"�/�a�%���v��C����G��,;�B�P����mx ����f�܉؀�}�l������8'�"���
S�R�p�p�-}�s�� '�9��BCH6�q��?�H�܄�þ�`DN�愻2����I��%5��(��{]���1k�J�g8�
��ͤٽn�.�i�pD�l�/h�*\W��π�����2�ɢS~�qsu�)�v�u��\�F�ׇ�.��֔T
�a�_���UⱣ�$���IF�W�2���B��Gq�&��|}�m��1��[~w6-�K���k.� �B�t0k�P�T�Jj|A��g����r��`��tp�� u��p�e$���Q��ϭ%�:�x��J�0�?L6ؓj@ћ;����l��.�G�y|i	P�v�`edd.��+����^���eր�-ݳ���D�%je\�����ݑ�H9� T��_�a�y�dHQW�u[gK=U���������>
.���Gcz{����N2���m�r���"�ΰ�'����
��w���ԥ���ȋ�{<�-�r�Th����[�>
%w?tQ�e{� �&y, �'D S"7E�&M���@�v��L-Apf��y���]��M�ϲm���Σ�@1��!r�ͪ|g��4ÆP���$�A$@w</k�8:U<���i~�Ȅ�Ђgka�2&�C�)�k���%fh��nn�d�J��f[w���B�N����C�*ZyY}+�Q�k�fa�R l&����:Kc7��Y	�*�NSP[���	�b��;����Wu$�B���&�;_R>���-I�/%d���_�C~�%h|��$�Œ��.�
gX�z�"�E�|��� ��6��a��,f��1A3[���Z+_/1��C�����a�ߟ�Y��_�T��	��B_##υ��gA�)�~p�d�(�~-�)􋆀
2�Kt�v�tyv L�6O���:�ȝ1R�"=z�D��p���m�i�*�H��0s�#P ��Ď��Ha��F�?%*P|��t�R��|���d��O2m��D���ʰ�t�Iw�����i�(�h2jD[i��d�ԏ�a���e`�����kJ4�j������Z��������}����QZ��8!�7��Q���BD����{��*�`2�
���ƙ�_9ڙ�Ѝ�7N���9���wq�UA:�.K�S9��Y�=�F�N�r��t���"k܎՛;�U�P�� zEg����?�|P��^7�ջ�6faTR�-�h�?��w��h	�#��M@p	!&���9�Β���ǧr� VG�_�+���h�u!GX��u1��W\.R���}��h��Ĉ	�;�Bڻ׽�r+��]�b��Ŏ�j��ݧ�u�)�DZ x׵�D���9ʣ�T9��V��,��Z�}�8
�����,䱜��LH�P&�'�Iø ���u�%�����l��N̵�%��dM�;6�1� �R��y������󸭺@�,��56�!N��RT�����ǸC�kB����'KO�����X��pijH`��OW�7u��A��4a���1~+�����-��Q�^�/
�=eK��/m���%C��<��k阏�b�1ˁ
C����%h��M�]�
/+��M���k�h��J̚V �x&�DQA�����G�O�t��/Z41���j/g�5XO��t4ur����v;�ũ�a�H����:����p�L]O�������[���zU8��b���3����{�1A�M9[��~$�:J��Ub!��_�3I���u����~?����9�s/�Ngꗔ��⼥�їl�����Y �Q�/ 6����/��y����o���0} @�G����U�F*�H;4P77�II�@��ׅf+>Eߣ�&�hBs�T���X7,�7�7K����u���jt4��#uV�nmn�T��(�?�,;�.n'��b��ޡG��w�*��5z(����0Yj����݃q�M�����V���of~,!9�$��=�3r��h_"`�'�����y���#1�9�����NP�	\+g%�n�����V�KM�<k^�i5�k�IUkV�ҝ.��bK�vb+ܖ����Czw	�@�~b����q����-�0����Q5�xބd���ZW& �/:֪O���Z�����ǫ�^a�<�*���g<Y$�F!����6�oo��n[��&���z�Ңՙ/O���A䴦�r�j��U+�YF@����%���}��A(�t�Š"mDs�.B��?����q��'�gX�iK���ѰdU�|�ۻ/�RX(�I��a�$�ݭ�R��x(*k2���"�5=�?WK3��4:�Ax ���o���lV�"��T�2o�n����1.F\�R����Z�fw�z��,(�~���v�[���%BK8�d�qQ����
[�5�\|�"ܺ����Xq���_[��.��k�ZY>g�ʅ�G��(9�g*Zơ�w��f2�A��K���*�F}l5������X&>Üւ�KWǔm=$�bv������txU�?/�v�?F��@ޝB�|�X�.��\�.�cD���3��B�H�z{�8��)�#�YjŴC��(�q�.���W*�UPֆ��B�lM��I�����z<29{D��!X�zz���j?4�[`T@Nˈ��xX���v�
�� .I#=i����{�Z5�v}ͤ���	J�?G�K��Ub�]���a�^fT4��,��AĚ�z$����k9����Qq0�����j���SIK<��"�R�d�����\x��	����ʰ-�N�H7�C����ߪ P��욦�������b+X@%�=�Z���_�cS�뀰VO���r@��X�+P{Vd�����I����&kJ�B�p/�`��L�K(�� �&�mQh�in�M| ����jH�DﴞM�Sc�/غ�����h���6��/�������2՜�B%�0�*�)T�O!�<���Y�(�ӵl�+����	���
3�nL,���2a�_P+6
���D��y̋-%�T\Y��9�U�g3\[0��H3�����ca���|}`l���܁��K�YƧ����.�P�w����9;L������@�S�������RjiS6�n���y噚sE��{._ϊPKL׋�Zس�m_XE\fGn��0�Ϭw� rW����]�{��v�C�1V�=|�C�%+i0����7hoe�oewu�g2�XxxV�����}!���"r1ҵӝr�L����}p���/,��/�kV�/7O����7�!�:�iV��^Q3a�n���#%���� b!��Hҋ@��ܜ�u�!6�P��zoDH���F�C��:���kn�$�F�J�h�6�k4%P�Ð�D��_��0�6F��P&��&X|�R�z�˨����ri���{���uL[�͛Ϗ��^&���`F��e�N/9J���jQ�z�x��'>����6X�>���^e��������Z�Bl��EO4��p�ɞ��h��%\p��x�K[D�ZƂ�(ӁL�*i�-={�ѕ@pX��գG0�����蚑1��u#QP�q��[-�G�k��h�A�ό&6q��pI�R9�B�]�y��ͅ#�+e��/0Of��)CdU6}=�5����?�V��jt��$H���8�t<��:��g�.�p(��)�]�C�#a!��}��P��`.��B�O�� ��YJ��|�#�E�ȭ5l`�A�91/[�.�R'�ݨg�Y]��}��U�.C����H�(M�+�~3O%��=!|��@��4�s[�`4@��4t�h[8Q�'��w�uE�y���2V�Q����I�"S�y�V׊V�]�/`ɲ����tuɜ���b���7��Iu߯�Ĕ�p&7��u��X�x�n>�[t=c���08scv��]���gS]�}��=tK��K�E�J���:���r����)��N[ �H���O���{��n�eAt�
(� ������O$�I���W��R>;H��,�$j��V�+�w�BJ��fPCy{g�k��;
�}��j�d�y�E�ХB���E5\�%Ĥ&��p�6(ɭ�vY�|�6X��ͯmE�S�\�`[�J?�j3qq�"|�|�]\ᖷe����)���&s��4VV؇h2�՜{�?�����Ŏ�T�y&�S�ˢ:c����]K��=l!�(s&D��v_N8o�,�9iC�:�s��Y&�b����n;BB�).4��
�GTD��BSg�Į�D����ˉ�q���_^�����D�4�"���%�ߛ��kX�E�j�|~r��T�Ʋ��J���L�:�c�~S�gR��aC����@�la�M*�o��
���,yY���m�hm�bh���D�Y�MM�=GCaX[�qP���BS�mZ�8��Z��C���(UD BL�h9�O��'*=�:�D��ӎeMh ��׭�Q=-
D����A��3��ƫ,I�a���7["t�Mޙ4�B�+#����x(ʔ_Z)�Wd\�zZ$)�_�<�A�,����/��6�K����qjg�?�{��8_�w���P��v���fb}���DsB���<��%39��H��H%�!y%���M9o���
�,��S��-��O<�plIe����,����b�}��Wk���5��.5tצ��H�������PJS����>�+n���1�{�;����v�B�������n�P�N�Q��r"�o���LHˤ6�U�a�5G�M%*��?��^��|	.�e&�{
���"��c"̩2����uS�!@�a��ې���(��i*(.@ꀕ./�;�N����d,=��H���:�?��;��C<�Dc��{�����ȸ\���MOm��`��k��Tٜ����;B�C�$��4��.�]P���5̄�*^��<�b�j���ÜY2s��2m������m���"�.1!`ֶ���8��*�����)ցᦌ\FZ>ąh���p�O d`.+������>3�C�l��ǡL:4��2vｷ��7�����1_�����?�2]ĉ a1�i9/7wo�%���H��`�2d���WQ�27�Dw��g��H� ����"�	"�A-X.��l���}����C�Fdf穟w�����VE�%RE^��>s��'NHo� ֬UF|@���ON*���d{�q�T�(�y\!^��7�9Ⲡ��JYmTg�µ��r��F#}?�� �J�0�$�f!��`/�M"�&+E�&��.��f[q@V����9��*!Pnb�s;�K��f⟄a��ߛC|1���~���\�}E���@���[`����`��c�"����9H���ų�Y´U����0w�/��L�m$�;!�SaZ�fa8�5"�;h�F{��%�Zn��7f��Fe���.���(��e�_�n��Y����#�����М ���NK�3r�↖���ݐ�H��V͞�x�Ο��ɉ�Z8�����Ge��|��&�ո�#o�Qχ����3�����!w19:�'�����Cz��|�׻x/;��_�t_u�mU�9�'N�wvhc����T�cP�j��\R��#�\��!�>;��G"�h+]�[���B9��6��&�L���&��!�Ɩ�H#`2�K�MtU�H�|���ǢT�~���_�ٽ��Z���xux�ɇ/��(k'� ͉4<.�U���V  ɾ�,2#0�Nǿ)RR=9�� @'��_x8P��
�O�R!;�Hė`�x'eOTǲ�7�r%����8�]�EI��ϴN�����;Sw���d7=�G'5>3�񷟡P�@	��A�T�r���NP=��mi,��z�⸖�����i��� �uοd�´kK�{���&�^ �����t1���.���SM�ڜ�!�'�:/��ҸJRֻ��� ��l��z�kwL�s���{�قY&���'�ӳZ��`�pQ����.������t/[3>�bi�q��{��t�)O���jފ ��iW-=�ʓ���=��+0�$����m�aa�.�Ӑ}@���� #��)���&9L�[���T'E�x�N.�޸Bg�9�R6̔FB[��y��C7�[��1�Z�f�@�t���9����./�4��ʎh-#�w\oI�M��$7x�����S�6���4�o��:"�>��?�d����]�N �Z+�p��#��[h�G��)fN��$MgNQ�ϵ�7��RS����o���(�� ��-o����5��d�B��E�9y�CƬ����X�m\�sC�fw�+��@1�X���Ȫ(�����lp�FxIm}y6�|t,]��M��?�^"���vz����Ѿ�:�jq꘏��SL����d,���`Ĵ%p�L� נ��jg��i���B,��U�R��BY��Z�}�����ג����MԦT��Ԑ�w9��7���Di@j�0 S#7��;�A��c�W��������G���^�k��]<ؠ��H��;�q��SZ��Ihߤ�](�ߢz��;W�"��q��m^�	$�)U��J��g�.-Oc_0�m �͚���yWF��4�����.�-\�J�r�79����@y;V��a��'�ᑃl���E��a��I5@}�Zt2.ê/,��_L�<�Z�08`��5�l�kc�8��k��6��<����z��S��QH4_�O�c3F���kBP��������Ir�r�tIS�9��Fױ��W��>�\T�X@�`�Jv���KF-S��˘%W9]�1��P�喙�M5*
wn�"�F�ݑ4����_vt��|�6�l˞&hZOY��W�8)J:[�i�o�TMқ�*��7���18�gc�^2��	��Y���K�bW�hb��[�pa0H����1��ZR�+z�vޟ�e�3�v?����~4������[���j��+`�j�!�4I*���+�@D2����C�Nc�����L@���<C?O	I���n)\R]�$��>�.�q|&@]ַC�G4�>�h�15����
�@N�R~����>�s��&J���'@�g�A|�.�.�F��,&���7��L׬���̰��B"�#?����dS�=����H��Ŵ*�F8j�p�":�G�:��B�Y��HH�����/�0�uBi���f=v~�eN{~�;��u�3��\��y���^�����f�y ئ�GL⩝�p0�~�#Qld�z�G<~����`���@��@�\�'��ٌ8� ??�����xh<���uO��20KT�ݷ̨52*I��F.D�Ă�@4�q�b�
�-P���������۽��ՊY$��@���� �ʥp�DF�g���߈>�"1���?��kFE<�E
0�����D�������t2�ә��ǉ�?��yw������Q"[�����i%���ށR��uW���[ m�%]�y&�\��Q��*~��T����QH=�y�#,f����'��k�� ���-��K�g� ��e��E񎳧�b�߄B�NQ;��S���t��[V�c���	�0� ?j'Z��v��L�%�$Q���'�"q���~�3tN�`�`�ͳ�i���cc  ɏ�i�ϳ`#X��m�I&S�O�&��H�1�v�v��p[Ie{mꟴޝm�;$(d�<�|1G�[�-�P��bU�j�4SZk�<�}�ځ����2c�9M����D�t�g]�N�S�8���J0
D?��Wq�܋S�D8��y��*C�#���} I[T��gA&�颜�Jc̫P �
d���q�o����&W� dp�#W�xp�nC�,�͋��A�l)�XU�˷����r�kBa�δ��2�ˇ��á������ Fy�NR�����m:M�7�d��Ĩqp��'jn)�����&Oُ��ɑ�s���nX�Y7z� ݈^���q^�Tp ��^���211q01NQv2�	������"���9��U�w�Uu��bÃ�ۂ�ܓ�.L�ƺ/F�����3�^�q's̥3g)0h�/?�U��O�"=
d8z5�@��3���mqu��̴����H�2�|��и|�=�tضj�2M�I� H	Ps����f��C�󓾠�ʆV�����+�K�'r��WL���b�x���d � w^\���Ԁ%	�!�NK���)o��/]�?��"��W@�3��_�o�1�v����!f�K�&evh��g|U��46�4p&P�z2���L�\p�9��I �R>��آ�7�A�V�^��Fyg��E-�g#�K�����HLn�l�S���}�΀Te�w��/��XjtQ���N�%�L9����=��q+K��8ߵ�ķ{T��ޒ1�
���!��b*���[�Ml�7�C_����nƍ�!j��d��UϛzkSr�a��e���߁�p>9�9�Tv��k�U���	6=��7��~��7ś�Ԟ��ꇢ��a�C���N�g�ka>�4u`��.���c�ډ�ߨ�&#�����˵��o�c�����)��xK�t?�;��t��JC��l�VY�^�d�ZsT���gAO���_J!���L�fpF��+���C=MI͉*�x�gr�n�u�9K��~�;�pM#�؏w4�Ա���P�y��h��A�u�Z���VNRCB �/�]j��D�E�{��������}ǣv�V�A���ݦ�A���	��R����WIb�xwf�?�+�Vz@��>�]������S�I]��0+Z��N)m�*��*7��4>�9�Z�^c�l"X�U������sӠ������Y���l���������éE��	���
({Q(W�Z�&��9���yR!�7;I�m��A);=6����G?a�I;�~�S.�}EV��ǩ.d���sp���b�O�Z�Ѽ�pg�L�� rk�2"��R�/�ODhF\a�1�������{1 ��� mpՀ�����*�J�B�*0W"��@~%I~��9��<��U�Ymt �ì��2�q���� -ه�@`^m���0�H�Fun�o����O��N>g͢#�1����)���k�qIi�6�g.
�����y�o�+Z홹V�7��F�������Zs�����b�5,ț~\�w��a�}�K�eM�K��M�Ғ��d��9�8��D�Ϥ)�>z�o�2D<�]9Ha��C�E�T�����Fvk�gI��m�K��I)����0lE9Vv_U6@����v;��oA�J_�}�x��[���6�5�\--��6v�'�y�*`�#?~�V��麳������?�<dI�Ώ��� Qͳ'�����~NE�6�?FJ��A=�7T,ލ�V���v_���r�$�#!���.���la꽶��� �¯����F:}C�����HUSs���t��_4���Y�Nf�4��ђ}�q�h�$j_sS�9^��Rtg�p�s^.��υ�݄����P�:~��[�n�՞RzOJ��M@kI�*��y\�ۮ��U�c�a���ZBc���Q�nw�jy�k���(��a�����M���*#2��$��U�O�<r�r�nFGĤ��-^ײ�y������GfZ�1ós��4��5�a��^���@�b4�U���3s���B���U�k�-:�s�)�-�^�+�xW�B��b%e/�����i�����)�P@(�N.V�Q_�v�!��e�#�oӃ�`�n�= .5q�:&�%����=���:޲"��!�软�\������x�G�_���ᇋF&ٲjU�Ǆ���^�,��~�������']+�b��Pbj���Ow�%Z�|'U��';�Z�*�\�R�Ul��EM�x;���m4�����`#U+O'U%�\&m�J�=̻H 
P�ȑ���+K�t�Fz1���^%��z/� ����M�e9>�[/AZ҉ȱ: ��bD�5�0@=P��$���p���8j��S�n^�v�E:]CXp��.w�� �43�}����d,��ݨ{�e�=�ڧ+�����m"wr��iiq	������[�嗢9t��~o��+���Ƥ�W�-o����,2��+}<�A6����2�r��C2c<Ų�h�ɂKh�/ͤ�%ଧm� ����p��(��v��2&J�P����ױ�]�!VMR�%K�o�R�H�����&<݋� Bi�[Ӎ�צF�U�4��lF>����$�]������l�{�Z����pkDN��q��J-I+y#0!�N���xBW���9qP�|Y}�]��ky���R���At�
H��'��Q�������D����s�a��req�/�W��3O0�d���w�,+.L=v�Xѹ��$�ƕz `�f1��Oy8���#���#⊝�8���+�ƽ�X�2TI������6@#��;�,[L<\�l����u��\��&Wxr���V�)`z!��,��xOjӲ1Z��]�p���C�]O�z�~KH���7���Y�m|c�[,���LIA�P�n����f���}nL4Y�hx6}�j���v��<��U������ݻ��2*
l�Cr�ip7� ���\Q9F��Bo�L@�,�q���"�!�(
�� �y�.��R�N�ID��y���z�ں+��h����E�8$)�)�B\r�M�vݸ2 ���
�sup&+�L8I��V��;�B֡}hxd,�������R��s�^a?��NE�u�ܓ���7�Ȍ��
l�t��Hcz~��;��C�q��YF�r���s �_p?�A�U�����Rv����i�6�7Tr+G}Y�Q�}�\CD��=���*�c��A�$|�:������:�u��U{�l�h��.C�Z k�t		�.����4�W��+!���0Yp�vA�ԥj$}�Oﯬ(˃����hq�����V3=wk�.U�ɃV��Z�ކ��d�ɨ �B3�->�Z�" ���z�1�xC�/�����:���.IoTH�s�F�n�DbK��ON3�1��:�e��
��"�w����Ao|;�� �o�Y�O�©�N����'3��^�v����y}�[�x�_�+���.7�� �L@���9^���)�F�U/S�<g��ZgD�%0 "�me����d���pa��@ed�!B�i�P���Jث�)M���Q���LSj���eW���DȎo�n�U�~�ْ�������G�
�R�i���YݷT�Q�6��<��=����m���}�����D����1S�e6r��8[�Q�����t�pl�},d�"08OD���g�����7Ys���eF2 �J�ς�M�:�����x�W!l3�_�ƽ�2�ߑ��i��D��#v��K6�<���ʥN#k�Y��6��d8ןhb:f�f��Y�]|
�nV�&G��}@�x�ӯ����&[��#�?�6�E��4,C	�|��0��9L,J�Z&1��x��.��:�S�H��8x�}��'8�����B��k�Z����p���f;�i����"tQ]~Ԃ�j�P�/�8�궸�������j;��o'R#����o������"${�݌�$ClR���'�
�d�hw����E{B�*���������|(x�F\����edES��B�����ì�&���iC@�4�m'���5W���Y|Ɲ��h�%w\�ƿdpu�1� \����?�Yes�=��P��>��0¥��@�"�d�>�a*L^�Q�%�Y� A/�v/�h�����Y�x�~� 6V�K��Vg�%�R�?X����(�,"�H�9
��� N���o�Տ��6uOIST�d� ��XCg�=�u�(k�m�<W�r�Ã�}����y�p@�f�y�T;w�T�K����:��Wa��S��xW~�1��w7��zzA9ALӤ�97ܗ����'.7���_Iwu][~�۩:I�P�ąH"����{X�R��h�?=�f�sH�I\Z�{=�]9t�e-�,�Vhi�H6��#��9�w�T�ao���sE~ܭЧM�����s��ܺS9�<E��9o�Q��Qy��_W t8��GҘ�1���Y���f6=��0C�f��*v&�Y��h/wO�p��	>÷�����ЫOۊ�Յ�K����_���*E�G*ˌ8@�
ɭc�-Al9t5�-�Ĭ1�fR���+L/� sG��{� }n������T�/(�e�6�_4R�:����쩑;�U��d��ה��}BT�hr�7VLkԊ*9w !��+!�Ƀ����U]�z`�P�����L���"�佷�G6H(��RЎN�<j���/�\�# 3�f����L+��4���(�
}}��bq�ݞ+�L�tC��I���l��c��<�Hu}_�li�"�ir|��z����e)��#�Lzh��?\����Y( ض2A��������э��Z���<�������f�^.���;(�@�<vI�Z�3<9��%������� ��Y�&߰d����C{�X$m��~�<N�aS!;ઞ�v���<���\RЩ��=� �c^�?+�#�ۧ����V����k ��}vAo^>�u)딿�RM�d 8Τ��e�
#2����5�o�7��,��0��L�R1:yW������Q���<�a�b��g �-闽ObykLRw�Q�\��n�:.�u-b�V��L&ғ�ٍ.��.�Qzƿ-G����2/5�W�ړ������]5�XR��e�= �~�JZ���9ߣNUUxI���9��'j ^JEP�d͇vJ��k���K�Վ}}��٩�����)A����W�V��i��Au�qC�Pd��_��s'|�ږ�>}t��Oc$Q�s���q��(�	F�EGr֔|����]t�Āt�����?U� ��%�Ҫ�E|���39����XU㸟�Q�ڱm]'�<����~}���#N�F}1q�ֿl�0��Dg�QJ�^�ڞ�%ؿ��j~D~d2(:��E%%~��TW���exO�*����)�ۂ)���1ز0�i����#U�zS"Bn<p��a9��B�|��崒�-ӳ� ���.Ce�Mꥄ������F.�زwD�v{�r�sT6�eg���2�t> 'PYܴ}1-�����DX쒳�l�/�Ǝ�o�'x2-&<:� ���`���d͹騺��g)5,� �5�-�Z���sz�n�p���ϔ,P�R[�E�A�s�pQ	=�ܮ"0?���U�	b�47�	�$ؖ�r)z�Y��@����Eqd��xD%�����^��J׽{���OܰRB�V,H�Ɇ�Nm��HjY Fj=Hz�k��&a˳N
�::؜p'�~H ZF��[��[�S@
L���?eH�s��NNGؿ�ĉu��Ŀ)���뽶,�W:�D*;�b/->�H�_��߀9�0�6k�����e����&��cn�͍���!�л��%�i��I�t���p9�7W�/���x.E(?x,ft2�y)ȣ�{VGz�^[ xO�+\�u?=~Zb��&/K����R�,�x
4��%�M��Ɨۇ\�1C �(��K�*hk�}N�煸3���JWT����!�Pa�0���?q5	k{�f�^*9���@
�e���Mϵr�����'u��~�׀b�� \��і����&�� �"�T������J��G`�
f���{VmP��CX�n�����3)VM���X�"'�Z4Lb0E�h������h��՟��!'�3��m8��r+|v���O~+�ccJs2��ܳ��īL٘pQ���s�߈�����c!pc���@@�+k�I��i��&{�=�\�V��1-���G�{�!e��Ƣcƚ����6������?��@qXJ�p�3�K��/1*�56h�.�^ ��������ט�eEI�{W #��َRI�2<�c�p�{���,�봛�$vKkk%��Z�Ëa\?�濯��(�� �Lt��1�o,Q��#�|�J�.1��������QJA��?�2�n�z��) A�+��z��ʱ�Q���q/!��.nmH#ӇJ���C�k,^q��\��������/���u�hm���=d\���(ǖ�l�4�D��3�9<���t�/I+B�W9�L�lh��1Yzb�-;��8^���<2�����{|��+0�uW`������E	��9:	��l�:x���֐��νk	xd u}p2��)!cc����a��9����/��;JJ�\(iUX�{��+�耟sec�诗��R��HQxnDˠ)Fv�B���Y�aX䎿���ح�5'��uT����g��'���|z����u��I�#�@������.�W%��N	�qZ9�����q�k�2k	p@�EǜP=m�Px�̪����<�n�y���V��:���
5fX5Yƚ\�ƽU�(=���Y�E,��P�����E%�V�	�ھ������4�c�b���L����~&�e:1���E��'����-Xz|�ǟ�3�����ۤ���r�������7"�F�w�j/��gj�h]���M���'����8�y�O~�����=��},���F-g��>ͺ�[<���R�;��ߌ�*� ��4��bl��h)���-�
�oX#fY���ܾ˯��&l/���9�:|��Wg2��1���!b�׬��r�\������(��/�?ƥ��EVرm�-U�� :� �/�2�Xe���%k���A!�d4�ɕ�#���8��'��}n-�'��S����aV8����i�f�������Qv������	)Yp����6[NJf9w年�@���]�ۼ6+��i���f�hh}��~eڟb	����ya~L�l�۳����^6�?�\�=�����d���0��<p��a�f��b��W�6\��+*���-C��.Q���������r�eߟ�m�:�tZ}wT.�	Q�)���L��]�_~�s��=��k���M�5�����0.cR.v�����ֽ�.�L��;��d�͠y0yf�O8+��Fi�W
U&�*;QM��i.���5���h�U(Q~��j(�Exj[J-ƌc��^4L�k.�tEM��oU��J/�^g����Ȫ.�?&��g���$�u����ࢇg�ܩ���� �����hR*�����$��L��y)fo�&�r/�
��Z�k���9p���s����h���5�y�H�ڬ�&�;�T����^WPg�����q(�߷M�2��|��]�A1���ͨ�9>&�q�ėt��]��Q�M��}�"莔p�|���/y󥶀��B�Ыl�;�����I����ؚ<%�2UI�5�J�ԋ����cp���t���E��G�)��U��yL�Vr �%�7ʖ�=�S>�P���;_blrz#�}�Q�	VQ�"�h�=_ `q�pK���;��)e����Z��-1r�d�V�'��D\�ڥ����"r�2�鑏�m@s PII���=�Ďs���6EKZ�?t�Q+�4����?U_����e�ނM�o~}���ܟ�8�cg3[M,�|����Ï�Nv�ݲ>���8�$����Ɂ)%����L��U+�ojg&^x{"\�swu~11�R
�KB��}�_@D��@���>�9ه�a��|ȲGY�C�b�t��&%�ut'���=��5-gY��"���9H@��ml�B�Q�ʲ�Dq!���*M�2Mp��ŏl�W{��������̉Ƶ�=q����m���?�8���1U�;b)��5����%^��8B�_�#_d��vTW%r-�3�Y:�W�7�\�0�Y6S9z�\&�-آ�t�f�BSʆޝ�e��)�H��:���t�����5�!	Vw�L�4X1e//���u�Ǿ_\ʋ�Xl��"��K�X�p��;��bk��r�n(�Bo�=~5��f��s91��N�ühd�}��1E]u<`t\��rDJ��-'�>���\�x��K��~z�)���Ҷ?��xj??b�2�'8���* �n��T��a���p���u�Z��4_m�Ԉ�Ƭpq�R}��{Űm�"�����{�7r�ɉWe{�|8Q�|���NS�<����z���v%�<)�k۲Q�����`Z���Wݘ��F��L�'D���{7Z\X� Aj�F	]��^Ɋ���#,1�����C]-�>a�O����1ܫ�ג����9d�uӱsͶ��8[�Eo���ϱ/���(�vU*\9l��^�M`k0�9����Ω��,��j�/T���b=��L�j�m��LD��HcD��]ss�ygث΁bYD�1�L���'G[r:.�>�p?
t�8~�QHJ� �Ӧ��ܒ��醞�WY��?Y�Va�lj!�:~̄�m�����&6Pb�Qę������=�5By���˂f�ˊ�ɩ��U.�v��PB��$�XT�{��肈8Oa�S�c��%��#cE��{$R�ko��[gd�e�M�m$|�L���l�vm:���u�=���O!8����jL����\� ��o�����Wu�2���4E�Q��v�>��I<P�],r+�e�BGI�ժ�z��;�
�E�t�����Χ��� S��J:a ]��X�M��X���W�N�d��X��;���IG�_�+x�DJ�'k�-�qY!g���֎�9�$�Y�C�f���Dp�&镄Ԑ��O~�W�ps�(f�qS:���CHdO1�O�\�$Fs�� �^���(����@�W�s��l8D mc�uM�Đ���{�ݼ�O������zSĔ>��4ם7��L�Wt) #h!�l��1����+3��*l�:�~�������P���5(�nCX�_�Ki�,{q�!L�fFc�K�^f���\ �	mR��Gk ���⇊ZΨJ�k�.O��x�r�6�~�-i�K?���ع�8ת"��A�N�>k�N�4/"�`^xh�zn>m�8W
2�33��X��m|S�>R	 }�uj�����47p�8S���t��A�yB�K�ŐL�p��5ȯ���F�j�4g�Y(�8*T����qhE�K'��9�NݞV��a6D2.\ F���Rv3�bj�un>.1�>��]���iZՋ{��!���_?iF��x\��U?�b�Fe�����*wnu�K�aj/A��h�]����6:�h���BhD����Y*�U��<\�C�5q�]'<JhdFĵ}�<p���~e��񥯊� l\3�?T��Ɋ�W�P���z��6�ǭ#���4�Ձ8�@E{�5���gz@���i0�Sؐ���0]ri\���KB�q�C�)��c��l.p�p�+%gPoz.�;��EO���o�x&R�������8W�,���ؼ�w�o�Q�{� !>�t:^s9���"��#��YٻB�Z�Zǉ�u����� �r���(�R<�����yq+?��-��+	O.���T���E���3�0�FO��Mr I�*���oK��P�/go?^(��k����Kæ��;~H����y�Y�=F�B�x5�RjTYJ����k/:�귫p��*LJy�!}��.�),/�)�2���=�$F�����y�hf�Ag�l��JN������~�A�<k���E&�	����ӳ�J<D�r��L�8�=��B��лf��]�6��v�5��W����Ʈ��v��h�0�g�<ק6�sK|��B��" ����7g�P�����
�1�uJPM���@��05k�,�ȶ�C�=�&�y��>�g)l��`�^��*M����#�N�f��]�a�kp(O9G��'�$���v;�*$ɱ�i����H��f����!`�K�j�3%��qغ諗��<dͅ�櫈A�͎}�Km{g`O������V��g�Wv��O1kW%@մ�t�m���w#��U��)_4�d�g���onv���i����c��:��q[D�Z��b�B�ˉ�+JA�4�|��-V�E�!�=e���_[/1ףuÕ�,4w�BX[�����K�T��Ia�
SG���b�a)��A�|��,����~	�b��-w�o���1���
	R)yՏ��^� NAS<�&N�:�6���+P˾�7�/�爠_�ނ��Jɨ��ٮ��-�0y�KSD��Uk��C?�̃�|ej��!�E{�f��E&�]���oZ���!G�����p�V�)�+_��p���6N��z��=�(^k��d�+�8&���V����d�%�ʅ�1����mno�7�`:o�Rsj���bI�<�e4�'����}���p�BV��'r�NW��P�8�2q&��X����em+.���W�(S�/5�m�t�YC5���
�RB�@��݋���#N�l�R
 �w�؃Mj6D7��6�σ������#���ZPŲ��p]�r��
�5;x.�#����|��Xє<S[�H�d:�~O�f�E&�{�s#��tKt�x*i��x�]�ՐC�odW��y��n=�^e�l/�ҕ7�hU���O*H>_�R38JIM���҆WX���vQiK=��ะ�8�����H��B��Q�I�k�od4������n[��|�$j
�HkR�@9�uV�'⼏'�_Nq�3���w��X#� eQf�婠�����/[����I�uz��`X �7��d��,��T�P)7��.r�/�����I���􌨷���	��;�<�%�V�$�����xG���=�|_+ϔ��U�%ݳ�ú�1B˨i���_�WU�s��O�� �vk�#���,S���[����a$�PB��|�pD��x���[��B��5���N����4�e�i��t�B�D�U�w��,شJ��A5�aي2�-M�vgK����X��S�xӊ��&�V��O���Ӌꃀ�!SV[�t�EZ��ԏ��t[�/�DM�;��,�;Pf����"YOAad��+hk�D�gq����R��YE�-��f]��JI淤���Bl��
qr��(,0��^+�@�Uhf](v��A��4m\�1�D���O���ybM�0�BM^4O6�T�����������LǘTuX%R=V��΍�gG�I�?�C��5��a�u���+��6���tw���p�J)��0a �NsD�9�8���<0.$�H~>ە�{%�jl�Q��Ľ�p2�PR:�����k�X�>zV�PkƧ����i^&��	�!;C�mU,Z����������G���o�}t���s:���%�]
|㉎�G��௞�����@��s?<1�6��QI�:�$D������A�G[�b?A�n�|���RELd��E٨�keO�6]��Y��X6F����F��.p��H��^���$��I'O���:���9���C�r�U�kᩓ%b���3Dl�����C���W<6 &��/��_B��%�$뿯�f\b8oL���95h�5�G�$�Y��p=t���ְ���M�M�����k�y M���Ʋe*?w0��L�#�^�S���~���2F�2�e��O#|���O���7�7��I�jiO��;^t)�B���=����2j��L�W�o�Q�r;����o$�.������0o�Pıx2-Qe�e��a�ޜ��lN����#H��X�bRݛ���T�&��J�R��p�7_n��Ŭ�˧���Y��M��,���F�X4�t�ɵ�V�~�p��,.�+�	�#��޷itƞp�x�jQp�\�ߡv�3��dkME��S�M�}�ʢ��"C������>J����d�$��
��I�A�|��1A�8�z>+�~-޵(��m�P����W�d�r�W��m&����#�2}��gN�l3J����O�I��Q������dP7p2SWz�-�	u�%�W8XbcU*r�9n�D�1�BG+�)yS`�����o��01Dm ~�e?E�'σ˽���UF�Qͫ�o�.V+�f;̷�z�\�]�������/"f=�$.�01�0�+u}
�5{�k��R��\�@�d�h�/Dv����X�,��p7#��,I�!��*�����<���zݯ���b�i`g=q�B���^}U���Ip7�i�;-��j A\�fz����|;@�ڞ8V���s� �_!��Q���?��z��;��<���[�Uh�W�1E�+��Lr#�㿦1<�ia�b'
�,�Y��[)dD��9m|1�R>�gIU�<5"R�����#Z�0�
�v�8�ɪ$�H�a�1��,�4>���) �b�������|�j��il��P;�H�W���V�J�� �:*��d�d�kd��c��c�����]\�T���ͽ�9%��w�0�;l�/��Ϧ�P��\5�+��έ���{12���Y����v<�0Ok1�%
�5�Q�� �Ɨ��7��Q0�)�U�3+��!
;G����	�އ��1��jp��6�Lz������`��Ŀǐ;  �n�{�Y�Lds�Wޝ�fGr����{*7@�[��=ZJO�JfǶ�u�I.�q��ɘA�<����"2��K�j"�O&O����H8�x���1�9��J��N���D���a���pFs"�&����ۅ�p����'V� X {��A;�G�jX�~�<�+� �6��@�["�},[o�ԥA����dֱ��ʲ���>��B��B��]2�{n��s��&,��.�`j��de� �G�`���t��u��ũ�Ȼ q�6�3�2��D��?5ۣÔf�H_�p%/1w��r�����c�|�3�1X!�6��G����
�""#�# �!�y䝯rf�����D�?�u?C��,��ߐ��2=�z#=�%��N��		���|	�vT�UȻ�ܷ��� �ϩ����QH]e����M9����R�ꔛ�m@��5���2���7,��d��S�nZL5w�kf�^����#y�?��9^��+�<.�v��}LI��Mwhʇ�L�Fa�5�tR?:�1���������4h�&�O��Rf�X�5#?NA�*���=t̫���~�=�x}?��(끣)�a��ЮQ�����߻�ƭ҇}7��^��Y�-�1XG�]��n���.3�уδYz��X���]�*aK�^S�m
޶�<�&+�oW�=�-Eύ�����^J��XE���8pH.c��ϰp'wb�֍H0;����5��}`����lMM��D��\SI�������z���>^�'�a�m`0n{�g�J�H�ҟF�,BB	H�~���\$v����YI��ձ�:��Y/��9�BX��͜�kh���\���+Jl�-���k���։�5�	�[�q��t�دs�Ch�&�ۏڇ�`F�k��sWt�r-�3����$vnU�Jp�^ՓWu�;8��/!���1M���f�N��^�6�Z��ÿ*30��$�ݞ��Z>�m��l��^�D\]�h&�rR���t�v�����J�����MPH4$Ў�>I�
��;�Ǖa�9�w���5�A��A�{k�-�u9�-R�g�,d?O}|QdA��NEU������>��>�I��R���z���%����P�="�I�[ZP��7����_i�tA2�[���9��;����Y���Go���絭b.�ɥ�����w��c�h�ssZ�9�W��嫷��ϣ�o�fF�c�J_��Fv��g��'���!VU��������P�侦j5�a���!��F�Q�[�yb��b�l�].	!�n��R(����4TC絃�p�tQ��RY��bW�6�����3����$8�eG�R4�h6�L�W�	���[0DT��Bo�E&=Z��*xb��5#ϼe�Oqu��6��aZ������.�Ck�P���3F�z|9#)�/��pX8f�ٻ��B�>��e6g�}���U��c���a���i}�,�7e�c!W+�(R�Ӏ�~�H��Ԑ}JU�Z�4�?˹��le��'�$�q��1�?$�D�.B��a�my��N��taN)�l�mbÌq���K�jw�,���i����b�b\>�9(Q��l�OhR9�nG�Z������(i�^��4���k�H�E��*�"q�b��_8A�<t�~]���s�!��R���UMv��X!�q���f;+���o�����
�܍�`{�RQ1ߜ|�P���u��T�J��o7��˲D��D!�g"��_oc~]L��P�O��a�F��7�`�����{j��C�8m�.��/���P3{-��$�'�("����U�P��5q5
qg���E5K�4sx<.��Î�.�;�V��@�nT�Cv�,�|N��>g���O�##��x����U}�A)���)$����WV=�_C�����J���&cK*zIR}ö�1Խ�'sK⣍LB�Cd9#�g6ŵ̨�'o���x�#����ؘGqo�H�Y��l�G��2$�zd� ,�qy��9�8:�8"#:��x�EIjk+8�����e�5GA��-��#`ث��8^�<G{0USO�/~�a礰/�x���;	-V���C��
,��/���C��-���&9jD@.�%2Km��r�COX�BzJ����3Bi:>>�fx��8�>}E��p��u<ki��m�2��ϿΉm[Ԭ������i�{���
Uͽ,��a��-����<5m�Q~�� ��mj��B���.'N�L�6?<t�H�=~K��g��P,�5 x(���Y�%�	��6T����_����y_S1���1�!?�i/�T���SY��X�H�
��_۪�����\�R"R $P�t/��r(��o�M�d����7P���ɜ�Qt�� 8�E�#҄�V<D�UL�)�0U>EY�E��m�l�����žAFˇ\�T�d����IPM!T҉
����j%�1�'n���2��ڍ��uN�����m�^���T�7-�sp�A���G���������Tai#�j�����wM�#��|Ǎ�_�h��L^e���1�]���F���<J�������̓F�~>;�G�fG9~v���E腨q##ą��>�h_#�G�
h�T��O���/f�4�����-V'��9���S?(io�����WtX%/'AJ1�Y��S�.:]>�c�t����Ц{�FKY�>�:���z��F�~]�`������_��Bʳf#p���ƫ�VX��5�¾��ޕ~�kt�5�ͻEH^��*(d��T>��5Ľ!�Nd8X(�\N���w�s�_���G�C�+5�Φзw���ahz��eh��8��Ō����f����~Π���kj�@���ˇ �A�����0[�v��#؊Y'��}d�	#��Ǐ5*/�JK��N�Wg�T4�VF�G�'/@d�w1*��qܐ.��V�t��zNw�Q"l{�ˤ����m��GnIr�����9�}kZ��Z�Y����_9��<�O���H'�5�����&�
��|w�S)_�i��h�ձ���
��^��CB�zp�~Ћ�3B �5��硴��3ӫ�EQ+��k|��u}x��Dۯ���h����z�z��o	��-\:��'�͓��4و��3����)^S1�렕 �(��ɯ~m�/Pe�d2���5��1�a�ym��b�r�3�>(���0��fs�>�T�2�W�1������KU�2����Y.�D��z�r#Yi�=l��ݝ'����%"^�{�5F���Bi�
@��="���N�G��l0��V��o�g�m�����V�zI�ƫd!B� �3qmb��2b+Fbwx` �x�0CTŇ�C�����b��2.��Q3K=503߀Gl�� s��o��#��]M�˾�C@ dYf$-��q�G@b��ц���5iˌ��{��c��&��5�o����4�)�n�?�L����dqyA��n���2�mӚ���	fu��κ�5�8]��z�|��붧�y�_��5�K�>�������͔��p�7�&^��W����o�!ʽA�᠛��Z����P�cv�HCY1v2��-�K�%�(�r��f�1��2���󏒋�y���O����tt�d��f&����⦷qo ��9A�\Yg�0v���_e��	���)�0ъ�u��㻗T�5t�2���[�>�F���QS�J��pNn%7:j�G��|��B~6;�����V�C��11Mf��~���i��I�2,�d��͊*:��>��7I���@�3ʘ�a#��^��co��2��/(���af۠r�@
T��.��`ZR7��1^`�V/C'�@^�H��������bP q}M�.��دR2�+��ڧ�ڙz��;!I#O ߿DSÎ�_�	=~��8�Φ��x�;'�jy�ϡ�����tiW�1��B^�L�]
Ԯ���W�Dp��{����*��o��	8��O ��&�Kp��ٶ�!R~�GN�8XuB��s� 7���q�M��f�������+m�XG���aFw����C�G`��4���/�ױ&՟)�\Bθ=�%���tb���|N��s|�o��;���m���WU�������nX�+�,��$g�}�eȼJY�_�䫱�d�zW1��~�M�.���N�3��%RE��>F!)^����y���]D<��_��>��6ZJ	xeUS[;�׵d�^�)����lLس��(6����f�-�4ðCu6;=���)�NN��Z���0��Ȯ Z#a&4����͛�������~l��t�����GC��5�a ^<]��{$�-y�}&��NF�O���+��i?�k��q��|�ȓu�5�W�~�Z�N��]'�o���ٜ� T�oM�X��Z?�k��Lk:�}��|��	_��qsVr�k��Z�G<��8�u���LNi��xU<d�m�m-�m �*�U�K��X1����������R	��]��NL��o��v��ϿY!�j&��.軍f�r�r�?�_�Z{�ý��v��*��-&q����EQ�Ch@XТ��]��!
�V�W'��5�Ͳ��$�DB���[��ZƔm.��@���2�q�ɖ��p���U�������vW�4�u:�tb��G*0@�1t�"<0C��$��j���'����<F�'Vt`��@I7bER��}g�ըFxW\����a��L�_�j�7��G��OWG��)ѭׂ��,&�\EBHZ��QR8	Oo��ľ����p�y�h����>ڠ4�۷}�)]gk`���x�A�`�1n�_REm*G �8w+�%�~	rڿ�J�]D2��5U,N+�n!�C�䷎����١������z5F���dC6�3�$�勖q�5�x��O��RѾRM���2�� r(�������
Rh1!�I��(r�F� ^`�t�Y�a����3[/('������H�nsy��]�V�eK�6%w�f�4yg���Ӆ���,2���Y��f�;�.Y��WFr�v�8���Y/���[����1�i�Pk0�=����KN9� �6'�����씿�R���N�{Lܾ[k,��(ʣ^��6��]2�a�k�W)��P�Osxa|���5V�c�����p૸L��$���Y�D�����,�z�-x��fXHW�|Z�7��zd����؂��!pT�b�+)V���3�ϭ&Z���F-�����ۣg���٢1�5��T1�F��j7��#M.�5@��O��@r�,|�?��˔a��e���J|cړ����x��Mj�N-��k�X+b�jx��B�l�a���Ϝ�M�v�ZJ�"P
���P�.d�E�=�x�Wf�<�Ep�;岉8�'H��g�����(S}'�Z}$c�a�*	�F�^�=:�o'�`Y!>U6x��@��vͯ1��ގI�{��d�Y
N��M���b^Fu���`����5��١Vb��F�>am\\����p/xL5����u�G׆;>Tn�)+�t�e��5�o��8ՄiTy�3ʠ�^�@�]�?��FT! ,�����O�S�H�Y��ȏ/w���ԏbt\f9k���K�JEn�
�=c|�� aR�Ej� DU��᭫�'1v7&�ռH�z�s�=-qiI�I���/�I΃�-�;A��.�dI*�#]Z��_(�3s��v�K�$��<���I�d�ї=+�Z�������ȕ�洿tDF|MLJ��=��O=V$��U��ft�jo���,�����nẽ�qN�'D������Z�	i.�Mz��>��
|c2%�&T�Y'�8� �`B���n"�����E��4�<��Hs��-�O0j/�1tāY75�TJ�M�CP���}��ҥ����xl�~\�^����GG ��w�e��U��^h{z�{;*�.!a�:�dTR���]��洶8҉�����fn�,�ޟ3 bIn�mx��yWo޻G-(h��<:'�c!��np,�#d�w3�k��`�z�>ɱA�I�2&,�T�s�a��+��?�H�1n��%����˸ؔ�īC�T�����������z�Y�p�ڬ��l�bH����!D�!Ҍh�s΋�c&��H}���D΁H7��!DC���[�+ ���d�5�UӸ����]�a�\�]6N7s]���79?cnwk��>�c:t��� �2��P_������π	Mł��cnu����/���Q�*:.��<f�v��G�5 P�4��E��
S�d�q��!��u��o2GY@�:���nN�mV9
Z�f�x:|��a/�!#F�EnǺBȮ���|Pv��"Kw��
 b"!Jᒘ������2��p)x�r�8P�L�X#�6�p�K{׽���i�,+�<�(bM�E���l�ժ��>|��%�|Y�%6�0��|,LܿF�W~��+�>�~���
ݜ�=)}��?t�Y��+�VWrTa�kW$�z�c��a�q�L=���m�U�V�J�E��b�������r�m��K��(���K�����	A��&����ߧD�Hh�/�T�����xk�s�|_�"����#6�*m���uTJx�+s�s#w�/�	���V�R��=��
g���wN��Q��i��(=�=2�|�3�bė u��A��|"��O.+�6���o� ��m�w���������Vb��gv�<�qh�'vQ̊�t�Rfl�H���4��7���~��a�̩f��2�ܴ��`��
tS׶�5S���YE�~wo����q�6�ĕ���J���z�t���M~�%���k"|�'��&&80�y�J�[��4�DJ\�E\�ݗ	di2�;#(�'P�fŤ��{U }C���f�)�6��ϖ�.I��-�@3�*�3o�Kzn��Z�gh�������g��%�7A-�a�A��h5�R+�P��O���bޓ��X��>�wV%b$dͳ�J�ٍݸ�P7įb���ĸ�.�xl���tHl��㙈P���2��tlΐy��h���
�!�f�[�xgMOR�"��;l�~1�k�<����
��Ol���b'�[͡^P�z�a)���\�L�f�D+�8.���� �7N��U��,��Y�X�T�����3��?�!���ׅ�w���YE�VR˲m �m���C����mJ�1،�I0�}�\�q83��0��fٰ} �r�lG��l�<Б�\���~�Q���^Y��/#lK�!��	l��Ѿ�=9�!��������Ɯ&�>aD�@�D�Z iC>�{�I�kh�$�uK���D��tP���m
`PB�w�|��ua��@�u�_/,��W�����T���QaՁ��2��z�1W�����&��B鴛����VY��<������/U��@ɞ�ᑐ>�8��w�u�BR{�e�$�67B+ȝ}��W��U�`�A�\!�Ds�@�uI/'��ڞG�a�T����mp>���72E�^��W�l�%�|n��3%���y��t!�u�6�.�X���B��:��,b�&H�h}����
+kp�q�_��.���7ڨ�xX{�x^ĎT!_V[�G�ZPW@��)Z�&��i�!�F��M�蚆�ϻM%�Z�
t���E*τ\���;�Q4�l�z��2[���a��/�m�5�_��%5�O���4A��A���ۊЕz��@XBCǧ�6���'�H�ϔ&��3	�p�눜�/K�z���8ɧ=������ġ�1q�EI���*��$w�͐�5�"J�+uDm������'s�
�ug����^D��M�	,(�zc�j~om Q�{$��}>�4R{:�#���@��g��&��n\À���Ŭ%��i�ֽuW��eQ��~��X\]J�"gK#�H����Ʃb��@����`�o��@�r1��G�#|�������
�>���َ����F��n���pq=g��g�T~e��RY bh�e	��񏜟�l��h�xqD���c�]��y8���3�3�y#�(�lf	�ͳ��O��n\�\�Ar���m_h���0�_Q��$��qC��J��=�]�m���5��9�(,_�-_�hhy4��_G�dҪ�NWr���E܄�Ҝ��Ÿ�⠮^�`*��v���~���=dp��8l��h/[����q�0����7=�L���E��	��3��#�7Z�����u� B�ED'S���`9������D��	�O�Πbs��4�#�"^l<>���돞<���Dl�i-/
�a�jc)��Kg�3�
�{�YM�X9��\��n�0x��\�Y6)`nҖ�^���%�a�ģ�I�R�I��4q]Ծ�Lg�[����!܍�$MM;s��"��(��pVli�����V:�x��e��i��B`���'��x�]�np)��P��Q��8sg�PL�}��G�4p�3�	��*͓��e��/3m�L��v���K�\��.�)���.Q�*ƍ��Gf�:��(:"����ѳ^���d_n��L��A2= >���w�K������8����ek(�]��7:-؂�i����.�jD!r!e�"��Ю1�9Z�$�뎁��&��Oh��Uk���ډ1����̖�Z!�,��3}�%��Dၠ=gs֯^���<��nE�b�����G��#nB���_n��
�YP�����k*d���bέ+ɹ邠��		}��`�U���v|猬E{�JevBZ��*�P����I��!3�|y������թaRc^6-�N������ف�\��3�#��2 V����P���,�~A.��év:�£�w��g���g���V�H5�٨Q�ড়�!�Φ�^Y��=A�|?EE�2�`Ь����@}7��Һ�T�hc�"�;�,��
`��R�k�u�m�#�1�d�"Eh��bp�&^��\uc�6"����|�\�����b�oE��FDk�e��	�� �w�a��۱���8���R#>��z����,�[�y+]/�[+@(�^�~�y����i_�|����@�	�)�Q�4M4u�Ӛ�)b^�:Y{�E��5y��،�L Aǵ��4'�e�f7Vj�s?y�K���gM��;�F7a�d�e���w��(�\L Ƭo�<��:�W1SY�<Y�B*^�y�839[���&i�|4t�GBd���`�vNvH,"pH�#�@��t�o��";ǥ^]�{�aӲlx�
��܂Juì�8����ȥy�N}���+�����{)��͑=ɗ*��G4\�N�BY�����.�9/��Eʸ�JJ�q��6W�^�B;[~{G�-�:	�&�/@�A8�Yѫ��3 (Dd��V867��D��w�kY����x�2�I�x����T1/�vk�Q^E������М�2=��D��J�~��G�GG�ǔ�J���1��.�i<��$�Q�m*�b�(��	����q2�w���j5���a��7��e=*a�j3%�s�&�#+�3�[~�I�BX�*��}	2�f*�>
'Чy�e�͞�,�i�3�X�m-L�k_�~��$���UH,#f��l��f�̦���8:rO�s����s�k']^�}��1qytx:jqإ�������R�M3�T�Z�e*�X$ݨ�(#^q�"+`>�4e�
\0[�8>��i�	��P֧��,��K��P��?$�ڡ�:��A��Q��g�3�G�e�V�ڧ��Z*Am�(��3���}M�;K�o����Z�����8��H��[�;	VqJ������V^�zKR��ҕ�/�[�+�?:�$6-�Μ��o˳�e"!Z8|�
�?�7�I��z���5"���o��+nĠ��׈�@>�c��x�;��'����<e���X��Tl�J�?�SI���1�>̿�m|���hx��f������v���v�8��[90�����B����f��A0/�I�t�������!����I���͕g�~rԒ����-�8`��e�+;��#Hx��� &��̏=9��]`qoW�*q<�ʃ=���R�r��'� &>�:+��\��(��4�%�q�;b�U����9����36$�W�F�����6j�+U���KT�9�6��s�rj�3;��i3�B!�g7�j�w?@Խ����$���\��aH&��:�8��@u9��������t
q1H��q�$)
�2�jT���I�O��� �(\S��������O_^4VKN�����v�}v��a{�H��mT�糝No_���{�`��J)?S�Փ�`w�?!��>=%P#�\���l���9ŏ����@x����Cb�/���i�Af�!d2F�n���N"d�:F�����RQC>��e �x�.p/#�P^�R��y�����n5�f)�P�\����_u\�@-p�CL�^Dh�O��d0^�5qe\�;g*��a(���@	n����룬����-�� �	�X���"�҂B��<��֒c��i�"G���k'�q>� ��D%M.��ߺ��)yg|R����ѷ��0��w�h��pU�uX��i�W^~��u�z�?�e�<Ѕ�a���%0�4�ȇؽ+j��V�&Ǘe��;[�,��!72/�7���kX�M5P��� g�^	"��\l�81�SN�u'w��]�/{��y$�}TMt1l�{9g/[�R���%�U��Z�ʸl1taw�S�ݠ���A2�AG�-���o?�Q�l�>���Լ�Ȫ��!2���V������=��/��{,U���]�hx%#-b�G���+�rm]U�J�?t����c�ԧ-N9m;�Yާ৕�C�T:.m�n���^W�VX�HT 	�lؓu���Eem��"� I9$�)`	�ݟ���힄����BФq��hR:�� /��(�z�y~��{ZP��Q�N�7��[�tV�b��Od�R��y
��3��G,���~�}F��.l���"���Q�䂌M�j 6�S������C�Y.���$ ��m'��!3M�����$V���mV�n(	��}Q�=��&y�喊�^r�h�r;/*��NR��Q��fR�&��;���~��YwtS�Ć�2+��)�����8�G�y��x��6}A������km�ZQGv��g��I����!Z��	K1�UwbHD�YCY:te�B��)W�����|���H�|�x �������7Ft����i���������Ա������T��m󫱕�*O~O&k��	#_����,h16o�l?�d�oJ�S>��)�t�Zl��E5���p���y\]��jD�>r2̼ڐ%�5���H?���D�#G�)OB��\x�ga�yφEA.�fB��G�	B�#��������0���E�}mqH-7i><��;ؑ�
D�Zۛ{��-��ϑ���@@�&�Ĩ�aj�x (�F�|�R}��඿�ُ�S�pn�%?��]���
L��[k�y?�f�J���~%����8�^���(����e�*R?�&�Q��S��1������c�h��G�jI��3)�f��{Ʌ�AM�&����������.�I������>Q�����z+�&
�l��a�t���Dh����A\ڶ�J��ã�^��39\�>S�b��C��ig��<{�M�K�k7���:1� �YT+�g�V�y���H?�۾S�?�Q��������e�:p��(��"����b�#��*���j��6B����S??�e�(�9�ж����h_:[aъ�,�x=��1��k1�<���5|f��)��u�6�*�����mMi������M�Q�������l��"�I����A�oV_����6�o	��� z�ƍ�6ǘ�Գ�����tЕ�<�����荭���ږ��Y6�M꧚%^0Q��;��⎖5U���Oc�=�2�L�-M�Xf��،�ed+&�%5n��Pm����:@��]����]`:���bY�'8̇?�$&-�J���TԎ�C~��D�PS|���xl,1�V���K�_�NI��C �?f�҄T�9�f����<��kSKj��|�W�n�A�㰲S��G;���j�N��np5�/ҝ�K�bQȞ䈸��LCTTT� {�s�\ 	�̞����p�0����̀ua߫���6�e��b�q�{n�<����T��+��Q7o�d�> ��C��M��pS~��\�dRN>��[�p�^�|�+�*�b����яf����S7Czd|$-u�Hւ]_����� ���O�JZ���l�E���~s�LĎ�wO�ǿ�Q�����Ʒ�|��al��1�y�MՒ�o=g3���[Ĵ��o����hG #����k,�����Zb��%���M����N�d�����Ni��^$1oY�Dmt���;Q�&��'8);��W��a��탩]���I(y#�G_���Q����m���iV��5r[��b�=��۳''?�>zT���
�]S.�\];�������t�4:�:U�X��J�U�
��iuV�=����1��Ȩ@�$���,���`#��� �����F+�!`�Z�F���M)E��G���T"V�܎Q�3][bKS=�_�����g��E �K.~U��|�rXѵ�a���6O�V`[%�8��O���f�TM��������j3�]���'U�_��F|}����x�߮����m�}�q���b�$�tXś5k:��G�y���l�gJ,��3Y����YyD]�Y���I�^ ��t��Y���M�J�C��O7|tU+;`���gu�Hf���вk�NaͣI즣��?Hp���ՠ�}�}��x,��L�ع�֝X��Ɯ���0~�(�^�~��΁6�Z�ֺ��}\G�%�pt�πv�<tM��VP��w|xd�-�[� v [�ld�n�E���#�3 ���q� ڐ}�
��* ���9�=�H	�W|�|��s4U�{���L̞3Ś�!�O�چ�>'�����n�:�6��gZ�g�6F�5<����a0{aFi'��|-�HG�UY��.F�X5�u�x�F̟"�������S�?hZM:}X�����dOK�����d�T�X�ݫ���ٚNП��∓o��t[%.�S����q�2��#����������W��Kd�YQ6�2[��'`��+C�G�������\6���i�p
�_��J;iW�˽���Zb�����(iAVƕe�
�shPq��()*w[�@���*�G�f���#� ��,)��g&:j������]�W���*>�J��6h���>��R3���k}�P��|����O��t)�Xw�C��Ф�K��E�OT��@O��EvDĻ|9iX�|��M��י��������\#X�~�_Q�������ǐ�e@LC�x=ۅ'���tX�w%@��-��h�gO��"�1pJ���ǄJr�9���6h(R���	�/�t?�>�,��2�4�=M{ټ��?T�8N|�@�� P���x�me�.i	�j�'��=?A>��ϸ��M�E(���T��hW� ��.�(kK/�8ཞ��R*�Yz:YQkr�7w���f3��]��ߖ���\�-s���g寨K���	��G�'="K���󕜈����*�u�V)�z����L�w�6�1hԞ{�Z�I�$0�j����I|���kduX���D��7�5��{q�9�<�ӯ����c.ɲ���?v#ĉC�Q�
l"T�@��ʧ��t~����@��*���?��Ť�
z'c��|�S6%O��M��W�y��P����O����f�\$�*B&����7!3�c������[x�Ue�&]K���ĥ�t�_3�Z���j�tE�Ax�(�alź�P���0�P�|2$�P����b�U��:�,ؠ��l6�qo���=S�M�����lOe��6w��(�H���U�۰W�Q-+'�5\�K���7؅��ޥm�#�v#��Z���жe���g�����a�$E~�y�2|0����������,��j[[
�؏�Փ:��RN�s���Zc�� H��0�N���߮�r����Nk3�^��p����>[�+����F,y�?^t����f��$��H���6h��9�қ��
x��&�x��� � �^��	ݽ���i���J@v(�����w� oh�n�J֒6_`VY�B�����6B��RP��UV��@�I��j]Q�M��^���lp�QЍ�.՚FP��j6��H�����h~�P��c��DUt�i���lD�G�3�r����_AF���C�����
��PRrftk�Nu��ia�I�����"��"@KλϽ�l��%C�d��ͭ����8��R��m%nL�{�?`�h!��ሏ�A"{���ƻ����f}�";}T�1I��=�Ф��;ͪg�Π�"�\�B8�~C���-8�F���7������^,WA�bQ�rO�2��SNGʍ_�����O���a^}%��>��*:��(@uc�~���b-�1�6�E�硡KZ�_~ �y�27�8	��O��l�`pa|g�C'���\�^d�1��;���lJ��a]ݥ�*z�կ�Kۯ�4���sMaF�M��)�8t���!�T}�� �PhpH��wN�;�x�A+@������4��gwH%)�l����ݛr����U�����R+Zc�7nFUB��|�71��/�ڔ󛶇l����i�Z�@U�+��:�g�sy/R����!��iK7q �:O�T��2b��x���zځ�pVu�&���H*�a�Nk�\�$u�s�k4�x��'m���w���F��ln�d�7�(�޺�Z}� 0��h��^{���U�#̩�^�Z[����b6/�[
�Đ��
�k$���ܮ�ċ������V���������P˨��3e����En�E�z^���)��8��8�D��#
��3�;��r��¼EtuX�*���%n >��'mW��?�ک���T�K�mZ���D�E����Լ��,&e<�qhûr�Ÿ��Gl�m��R<����$�b#{|���'	����@eg�'.�tߒ��:�}Z�'�C03Q��
����⍜B@7���z��� �y6�;���!���@�ۜ�:=�ܽ�S�닼��Y*�-�rLX�Vh�D�s-��!�0x��}�0���~p����|������ǜ[C�P�'Tfs�@�+JX�V��2*JB`��R��\���M�/��x���,��hiT�k�M	lkV]��=�8ot��}���[c��(A���'��Y�wYK���yd��솃��Y���U���OiaWJ7�L��d���\������#�B��`ܶz�����z-����~|8s��XMG��4%�VJ��*�H���畁2�2B`c[EO�>!'�bM� 7�*y�R�3��΂���ȵ "��vcp�x]$�6��B�|NN��l�4�P�t
��w*���{�Fx�4f�
Q�w�%��wDg���p�n�-6M}:�`�R�����`bU┄�'�ߧ8S�z�K/
��|oU�B�dJ��
\+m��N.A�`� ��2"ւi`��8��#�I�>����~��6�)4�&|�6�{��y�#�҆ 3Qx�m=D��0�,q���3�CQ�̯�A=����M�lM�˲z�b�3��->r��(O,�Ho�*V}? ���jӝ�C?�e�WJ���D��Ԭ�l0��NK�O��9ky��+3=. �K�}Lל������������oa����M8�F�����Cn*���"M�xzCXmsD�����֜��A�0*:���r��uz#t�t�M�����C�=�5����lUߗ��'��E�bj�Y��MxM|J�A	@(���TP�IDS��05;��^H��&C���d����j:��7'�>cEGR˾�C��؂�y��J�_�/��j�o�ê��۾Z	�b���89�}�k�B�V�KH�~"9(��W�7�	��a�?�����F�	������٨d��Ba����Ň���1�u�72��n4V����6���g�߆w]��l�Ru9ӏZv���@�K�Nd��
�@�,�Tex����'R��|:�,ԛf������Ei��׆ٯ%C��eF[֚n���a|I�5��ۂ�H,,�[���'8�۱��^�Ͻq��={Lzm���O��H��z�
�٦ǳ[v�+��٬��tFؤ
�9�L�2��R������ϡژ��!M����+��U�F<m_ҩ�޴j?���ٟF�����v�P4<�l>��a�W�O����#K+z
�K����/�����G��>?&�2��&�G�L���<aC4��2��WC����)A�"��s�Yb�7M� ��v#����V[W\^1>��a��!�/��F^�s��3��w�ԏ�93�`��g���]J-Kjr���s8� ��n5f+��<�ŀ.b�3H�<a*5]΄�k�&8�5�nȴ�P��H�G��5�\�u�E��`%����T�;�޴���X��,ʀ�|>q)۫z]T�f�`U��?˥m�t*�K�f��<���_�NW������q%�|���0�"�/%��$�T�埫�f��Q���A�^���Zo�=Y_P��C8[��q���}��F���D�3\�8O!�*��ީ8v��^������N��Dœ��$��`�:�O�]���@J�B��I�B ��.��aКU�7�f����F�?��Y���\���C;�����+5+��`>�)G�[���l�l�j���G��2~ٮ��pI��4)Ӂ���G��Y#���w��w��������^�����:�C���n�rs�L)t�$
<���]���ŀ��n_�{� �i���l�tuV|XL�Q�����Cdq�h���A�|���Dj���+�j^�a����@���\�pd�֒K��jox���|�=����]�УJ���)hrF;�&e%\k�����#�%����ƶn�0�祛G�OB�a�;Ɍ{0�j�>`d�^��e'Qp���q^y�y�� J�k�7���(���S-;l�%Щ�E���Pn��������.���W��Uw��ǔ��`�z��-�w�Dӆ�"��@94!.l1"-;���(]Wl��nn�Z!�>]�jW,�ԷW�d�H&��iH	�*�s.*T/2E�ᶄ�n�����f@�$a��@�(o�4�@Vx(��M��o �x����Ր�-u��}�L|�7�X�R�.l��;|Ԥ؋�	�I �h9PM�B��écyG�~���&��a��3wC�s�%7c��*>`Q]~�.�{���Y���}c�>�a�P�f"��-�>���rN�#tl�'p�婣k����ix�{s�YV}n��F�s�(k�y���MlP��=0���A��A{k.��h��^%R8�� T�wm"�N���%3�K�C�)]�in�ȝ��Ȕ�� BU^��*4�T�WM�Q��!j��rF����S*�_����� �WB�?�m���@�
10��(`�̟T#~��!���#�|+{V&H_������om;8��-�4��`~|���i��*�F�ӧ��!�v��,�a0�x'	i�����`F)���
?|Vt�ʭ��P��Q���T�pZ��ܪ�7�W��@�A�%O�8,0gDz:�E��B�)��
�������}��LC��&��<���6=�K����❢��
e�����[�!�{�Ž�̹ho'[�� �c!��}*K��&��Ê���z%��QEIO|��1m��#�SQںŨK��k^�VɎ�QZ�� ��A��v�L���Q�棪@(�y<PQq�]'e0������`q^�DyU��i:�4����
�G���Ԃ��q�V�p?"[����l��ӇCX�G�Y���0�m;_�(Xxޝ7nF0}�/J�R���4� ��˿Ώ�[|����9$�"������6��t��M���͞k�?-���6C�������:{�<-�e����Br�Ј옝����b�0��>(�{9�ϟ���C����X�x��-�Υ�ʺ�;	wZ�݆��;\v_o�B���@����	���z1�Կ�� �:<jl(����eB�M��r����b��G���r(�V�Q5�b�(�Y�����0	�G�FIk;K�<ݷ�)�=l�d�Lū��v�Ns6���q�bi����@��wz��WMr��3��x���0�ʉr�/��뭠Ű�|"��E3�Kl�+�/���O}���憆`Rڐ;/N��BB|���d�*���"
��X(����������.�e�y�KP�T�=@�$�c�����w�O�����ˠ�ig1���~� ;{���+Fo�%�}��:*�ƌ%}��3Ծ��XF�����̼��:hK:a,ƪ�E��&�իd��KA�����7~c�h�[Jݠc����V�J'�9��ZL�qq���Kví{v��W���q���)𠻙"��u�B�mOWUQfݢ�
$��{G`������p�%
G�(>-��$�n�(Z�e�r��l-r�c]J�`5��ee|����䥱-��C��A����-������[CL�}W�5u�}.�R��0�����E������N>Uj(�[���إ�ͦ�M�]R@Pg?O/��*�٤����&��7��FY�"�Qܞ~��ҩ@��gT�'7����jӏ�%���#�9x�B��2,�C�i��H�{��9���@���c�����p�q)�7~H�}&\8I����V�wH�TH9��XB�P�m��)/�y�گ8��/�k�-����
�h/�&��X*�(Hs9������L��1�Ld�3D=�Rv�������IST�VK�X{�r�B��e&���ϙ ��l;D�5`�>��w���w����+r�duo�!��Kg�����	2����4iH����N�g,�)�
L��!���=NdO��ړ!߽�$ʦ���P]�^f~qwN���~di֟�'I��\�7��u�@�7��K��}�w�<@�W����%s���NM���Q��dՏe6�3�H��Q�O�|��6LI��?Z�P�p1]Mu�}��6�hiT3ǞW��?z��A^yn޶���:�W$b�{܇Е��f�Q�^8:G�̈́S$����z�8��YW�U�~`OC����7�o�яE�y�r@2@�T��{��3�C���dqudE�`*�[�Rl�6���X5F:�xB� t֋��a����	?ݴ�i�o~��X�s1����X�ۆԠ�����}u �4����9ؠ�&�T�,05��`���)�� �Y��������W�`�G������T���A�vP>[�L�?�ǲ��>d��ʮ�ó�1�����t��1�U}��f柸W}�Qjh�٦����"��ʌ[�gTp�ěS����H��lH�ڱR��7��w�i0���:"�b=5߁�D5�� 񉑠V����$/�Ϸ�~�&�ퟠ��K<�
���	�����T�֞�-��4�a�_V�� <���-��L*53��d�n��+<Ȋ]���V�.,r���)�4��U;�0�� �!�b�y�j�V�Q�(l�-�.X���S& 2�N�	��J~a����̤������P23�D��L��V��tLs��f��ek4�d����� ��!�U��֯���ST+�oCޫ��>	ê���	���k���VZ�N���+�z:�*3?#�9l�Pykn˻/M�$�>�k]q��{ܟQ�wVo�ΥRWn()� ^�fޟ�~Z˂Q��)e{dX5���BL��Xc$�<�9�;�G��A�zh���.]���B��(i� ��S�� ���[�����9�i#����Jr�O�@�� ���<��C��!, �`��z%;|E<�E�V�9^H0�+�@��S�Yg�,�C�b�u�	4HX�~W��q��]^r�ɔ>�J�c��U��������%�W�8���<؉ZTǍ�O㕫K��apg0�J�[?h�}K�uC��2Grg�IS��{[��T�BaR���h(+�� 1�ٔ�@j���R�F\u�L_Кs�焣��
��b$�v�c�P�=Ka1_hE�L"�M�c:�E�cU�y
��K��2XN���� �8Wl�j�K#��u��T�}G��p HYjg���dW�s�;X�@�_�1;�5��j^B��C�f#�����̳v�;cq���t?'�i+��N�� Jq{{t|�I_mQ:l��af����N0��*�dR�ĲE���5�db�.�b-(:��L;��+u�`��sȹ�
�6L�_MVC�}:�T��+�J9�VK��������bE�Æ�l�6 �Q�؏
�UPYS1��>��P�+�)'����L��k�^�o0�!�]�{��\���X��7�N�@��nq�:�{?�L�E�H�r��@����(���8��4U�x�	`;-�t+쐔<3z���x�g�����A��6���g`���:���-y_��d�w��E�T��q��>Q}�G�����u��by���w��	j�M�Q��<�U�����wRjZ�΅�-F=���H��56� A�|�	H�Q��=���OSK6�?4���f�OA�>(�Qh��Ӷ	B���]ڹ�}���@�u#{Oj�Q1�t:���zZ�,�i��P]��bE�����U�e.��"4)�d�i����螰(��+n���
f�{�%�麧���R��4��ؓF6ط��Z]���K�	J�<�O��e5b[�Dmd\�6U��C<�X�/ h�hoo��v��!��Mb�`�2�����[�o�찭
f:�M���>t(˷]?2�P3�c��W!*�R	�0Q��80@��T����;Hj����V��4gJ]d�a���+�%!��2J��l G�Y��p���WQ:(X	�!�{.K����=�x.;�} ����{!��|0]PE��?M��b��K8.�����b���Y<y�s��?���z���2o���(@�~��A�x2�H�c�m�����9b4�c�y������#3�vJ�=�%�y�{=����\�� �A���C�lJ���*��/Sӭ��Ә� ���"����σ	���L�m�sʝ�����' M���~�-Rs�N�C}k�(�x��k_u�#C�h��_�@)(��+L6�zc
�aT�)����az�	!��̲��z�(8�O��,��t92d�����|[����&3w��Q1uW�sY{V3�~a�q rS��t��l�?�x�A�H���8���/c';i�a"��"0� �'���y���K��Q0Y��ū���Ο��*�%�(��$�#�S��Ƒ?cQ���LT��f�[��J�"�������:~O:��z��c���4V�Д��Ş���AJ2J�����K�샀��&g�/�ku[��Քn)��)���]�$���fƍL��N�/�@�KF��m�B�_Z�B�Nd�MB���*�E�J�$3M�'�S�Χ_^��xX��^��HU��zà0� ^�<���}��_�����ܞe�s���*�T�y���iC&8l{g��=�i��;�}_���9dP�Μ���_\1W�Y�ka.P�ɿ��Ks.#�_��$�6���l-�(C��U������ͪ�$5)MWR����b� /%=� mG�����X3?��TG�>#-eSRn	�:s�d�e��3�8$�a��;R�J��&͍RtѮ���l�%��q5�|}����FF�v{M�
5#`�
sX�|$h	����?b���_3���e��)N��M?�>�$��Q"�9��^g-9.ظ���-fp����kUSu���<�4�wc\����7�`�[t���Ax|I�l����n�O{.x?�3��A�紈5�=� 8��f��˳�B8��AXӖ�h�n~�>�n�#����+#�8�r�)O�Hꤋx��.��h����sN0}��,����v�������"߿J����Y:���"�2�w��?��$50�ջ���R͂�w";ߖ���t�ɫSd�N*P�Ǥ�_@����D��ٝs�G�!�aC�6j:��(Kv����*?��G���9 ss�ʢ�2@x�N�b�r͘bF�Gˎ���o�H����y̹�~C?��ӟk���[�Qp�>=��5ŝ��uv+BW@�f���:"�������`���݈��KM�cEY����Q�X%F��E~)�--N�껵g/�t�Õ��j�'@�p,%}�y
8�:������_���9)��|x�J��6r�^�Qz��8��������M=�(��߂�7)?�"�m9H���`�g�f�f���R�֖Kr�λ9�:z�U!�6�L�m	�l1���b7؛���?h4J�D5�Ig�l���	��2ږ�W6�u���*�1#}$�(1�[�k��X}&j�?s������?����f'���3�说y� I*��� v_;�@� "������3 �^���6.UԪPw'�u_P�+�+�ռUx��a����m(�C�����`R�S�H?�O�1.��3씐=ъ�0c�X��}�	}�|�V���꘲oH��HU�:��N�/lp��t@�A�;DJh_�ڼ]��L�"��}P"[m��W�X��@�ʼ�hT�Q%�Ǳc�@J?'��D���悏��5V�k�N�񖸺���r^$T�97=	1���O7�&�˃��u��K�wg�/_��!s�����2�y�!]�g�G�I�h�t���>O ���YqV���H�1h#䛠SWY��W�Hq�@���n;0*Pԧ^�a��������dI�v������RM�ʠ�=�i�X��J O� ٝ�AAc�F;a$��L?��?=S�o���dQ�����.��^>T�v��FqU�y�e��3j ������X���tm�t�Ih�s�?n�@U�ck�I�qOC証+�� �dhH���=�G�(�^���r��q4�I�v����Գ&̏E#(���fz8�F��Ue#ر�\I�B�UВ>�Ɨ��?P�F�/x�!q|K'cx���[-)�fcv��2쏦��`0���(�
�A���mq�4N�T��>&��@��Ɔ7���6x*��<$0�u�s�oo�(���r0)�]�J�=��[ΛD����gf�*�����w���Y������'6&���|��2��
�&V��"�#�["/��Ѵ����ݠr�*�[=Y_*nJ3�d�}��{1V��(R�x��Ԭ&ud0��,� � q�68Hu�m/�q������$g�`������	�h�-!c4o����ɦ��ԝ��n��5c�r7*�p)��=�Ac�J�7c��>��RMX�V�A:�x]W�|�7~½$�����z�V��Ӽ�����.�ЊC��G��a4]I< ޙ;�H�PJ��)��Te����Z��ʶg鱴���3�e����4lT�|h��:��o<*�_nS]��RIm���E\|�3�ٵ�c�M^SAGAR�����������^�������`wp)~w楻��Uj�x޺emc7.d -�`).dS���x�@߯�lM�S���<9�e��yI/�C{w������'�.���pc� �J?�߅�+��<g�͈tG�i�Δ!'D��	�2��8� j�6l�oR�[�G%���A�_�$O��P?6��>�٧@I��n4�1�N��C��LϿG�h�V��B�k۾��gW�~j-	q	Q����Z5 $������iN����8G��v1eNl��;�aUO�Z���,�T�0u���@�XY9q������!��ib�\�)L��RN�&��p����C/��J�o8��暭�,�9�C�=3�W�w�Z�t������K�;M����Z�q�׼����N�G�7������3C�{VT[X�r�2o��f�9l�dE�H�b����w��$��3�#�kKM፣}�u�HB�����2M����o��?���4,[�s�3J\FI�A5
J�����'�_	�A��x�܌3�����?H�2hM�I���Y�`��U��e16ݽ�>6���$�=�}�F|�m��W$f���zrP��T��>:gÅ�.f/�i�A��h��R(���ε�����
�uP��e�f�f���|���O�������W/�KK���)j�p�C2�E`�U�L-RKe�Q8�V�р?Ȑ��d�%M����4�X�v�@�%v���HK����^Z��Ѣ@�dD�u�_��z�����L��a�@����4��F|9�,>Ξ��`4{@&����G��>�C�u��6ʒ�Cu�$>io�:�\��`f���C�h��3p���W��y.Yx�'[[!͚x���v�n���D5@N��+�F���N��v��c#\jRu�wV�9�Qz&�/��&����
3�r���$����5���4=.�=��U����3�0m�i5X�/T��;��w����/x��q��;�x��A�I�yN�|��,*�^��q��Ng��Γ�/6�E|���o� #�J�A�5.� Ghi��:e�>�U�?ㄺ��,�L� Ѷ�[\)�����D����R����ܴ����J��p
ʴ��Gk%dh�QT���q*�ˣ7xN`(��<�=�~
�HVR�s	�ڧ8#[��8��srm�EBn8�79(�^��V_�k!?iu�˯��SX�i@���s���*M���o��ɝ��H�N�h���'�c.�8A��ǯ]�ݧ�4�qpm׉Y�Uh2]0
��y�u��)��+�K���BR���3�^u@2�ϲm)�Dx̍�-h�Sׁ�G�`&���b����NMW����5ϖ�j^�9���kz��ؚۛ��}���l�o�7���o�̛z���D%[,���LN]܎�S
D�T����4^�4�<��jh���F'p+�����G�FlkQ6N(�����eǖK�WgJf�m�X՜����t�����yB8y��	�"G�d���_kW��A�������MD����W��'e��K}���PD�!���Z���{��d�@ORo�2=?��C4y@(�΢��px�x�<���}����7!�3��3q��k܍W|A�'I|�=�݊3�؏,��ɵ���X�O7��M)��_R��r�Q�4'?�*�	�Tj�_��⌧��ׄ�����n,g�T$��Αֶ�!7�>�,LyŁ���'�/����B�;_��e�Ա��$T��C����i{W���I�	jU��Х��6Q:W�&uS��������SP�=?�n�>̛�!=˹*�����V�)�7%�o�V�UOn����]`�y66*jջxN����M�r�i��n�|+��^����W��de|'v��������ܗ��c���6��K�/�n����(��Z>��[���v5>��.���3�����p�_j���y��iY�P���-����8c�k�)�^H�g,���`�*�BF��5tN�;����H�B֜�F }jS�.�«Gj�|��K��)���5_PK�����'��[�p�S��[Z�in%�������.Y-6�# ��:J���nK�b�>�xߓ��P�@����!xف浲-��/ׂS'bS,6�0��3А���L����:y2�L�4߸�����!�ݡ���l�!�	�y���(I���
���2n}��Ey$0��26*AB�J?������o�~�h�z��0�EX�֨�!�*∫���m�V�Y'K��v_OU
���ǂ��Ov�}�}�n�o���Ǒ�Q"�	�a�����˞��u�����VX.�;Ċ������h�#���V�c:�q5mO$����H!?�%9�C�f:O�9�P&]-�ڱ?t��m?"9�qk�L�'�G��y^��8����;�yc,�������
5��.�낔�F�sΩlj)�/|��zC0kx!���n@��*���	��ۙ}�c���J��S>�0������v.��6��2��o���-�9�$�����:97Sa�b��ո�:�Pu���q�W;B������w3bE�ow���3�h��$�l�fA��g,�qJZL%��)u�����<3�·�Łe�̤��iO�z� ������0�@Z~E��E�js'�d*�M�\7�{���Ado��TxUS p���rIP��7m�_�AP������fȘ�������Ys^<�x�����:|
��(vI@���1!͘R�xM�iq(>e+ӶF�m��2��dv���=q� �;*��aA�,��$y�L����e�����=�;�����rw&���HSC:Fu}���7�v _@ӷgl۪����ҷO�+>[�U1tϑu�cԽ�Tv��Pr���8@���-��I��oh!�ubS��\���܇҅�BW�車qY� �����+�I.�L��<Ѯ��M��^�t4�nb��2�(nɠ`(�E*2'���k�H|F)+8R;��,�L�bų�>���c�����^�S�nh�W������?��4$�oN�r�о=�]��яQ�I桏C�7�]*�g���� ��ku}�Bf�2G�5__z��(\)��6�Q��tBu֣aRV�`d�S?C�R֣ՙn�p���J����@-�K�,qEs9�*���6���d��΅�Ki̼�W��Q�R�4uVі�}�w�z�M��X>�4�d�=�����>����cg����P�񏻫Tj r ��1z��o�E�ݦ�sVJDu1�C��ŧ)�����`ydN�T�s���]D�k6�5�(,;�@����?����ȿ�A�m���M��I�ړ�I�KG�_���)����C���:itX;]��^��$��{����@@���P������ɩ	�e�1H����� xǩþ����0QRi���+����k��>����Y�vm�o'���'W܀��h���ًT%;��y�t�'7.T��7�l�=��*��˅��;@�]�Aɤ(Z�f�~�RQ��ըt�/�j��M�
���&�*N�����3��ڊp���T�,���-bV�p�ݦ��kU�>;��	ay`�G�[
�W���ѾFq����7@�`��V$��i�k��Ћ�2�0�2@ ���|����Mz�\����(�y����</�c�� ����tY�@�����ɯ�z6޺��7�ʤ��"��_�cl9t���v�y���=�o/�_�Q�����<��D�6��tD��'�������ՄO����W�*s?��������;�.�W�6 �i�G�����.��:,��ynls<��J�
_/�������+t��n {�Q>M"v�vn:Ⱥc��+�jc�s��y 3~P�����$�ȱ;���H�蚸�"�xy��Z���X�,��1C�S��.��wΦ��[��g+�p���G"Fppņ��j{��<����x`���8Hx\U�:)�3�7�����R�}Q�+H�i��G��8jwƶk�/�S{�3�U�0Ŭ�i<U�iv(�9�[o�f��g=���4Ł
�M$�Jm@b�'_�!�q�.�ͷ�-��v}�S��t��.Ϩ{�5�b��$��BTK|~��_��une�X>xH@zw5�j�J"�m :P�w�L��n��^hlj^����P�῅AQ��A��O#���Ro\��Bo`�IGw�AJ?��(fQ2r��֍�tb�<��<M�	"��"0�.�>�d��}�O�_�\��IS�Cow�`�a���>���:�{l	���.��$���g̭��T���{�BS��{�L��E
�?�E�Yg:"�͕t]�ĸ4�Q����3 ���(WՆ��s��@�T��6 Q.�$z���zo=��i���#X�ý�%��e�1��>���gF!�ބ�%]qM��{ë#�M�,m|�>J����	�g�vk=L�����uCY�f`��4��6�ZZ�y�^i02��x'/��6�\;�z7�QM�9�`@�#�MzJ΂��x�f8�+�GX�7D���m����㾘𞭲���7�/�����xLW?�a#B�n��V�� �x6�'o�8�#7�=k-`�!*�M��\��I�~>c������@Is��4H� �/Υ�)��u�"�z%��.�_�^�]�ʹ�4N2�F���X>�_�.��^>`X��9�/��n"f�>w�Ȼ�f�w����U��֙�F���7g.�Y�=���y�L
I�)�),�i1󼭐�G��� X���C�!1�U2��v��D��"tV�$D�����I��:���;b*qI��`�m-�*�uT�λj|�/1Wo�ho�J���i��r�t��� R��<���#+���|b�p�,�d��jN-�����$]��!��U�Z���z���$ -���j`P���M���A���M(T�Mɕ�>s�է)K{��h���+)���cXe�k�9�fͫq��io7��	Eh�l1,G��bL+z��[C�q91�63�������B��m�&)�H����H���.,������\iu3���44�ӜX��?�Kk�O���2m�T��{�%�0i9�
�*�.|�)�B���H t��O&]9�����Le} Li�J�-��Dm?c�[n��kL]l�f1���_�C����R-�RQ^��68�x�Ծa�w��-ӷ(x���Q��c�s@*�P�����s�!31�c��"z�e��rt�?u)�yA�%~��a�~̨ұ���zZ�e��Z[�J�3N��+�S�Exn�?wU�ܟ��x�R��P�!B��4��bT)2Z��:睑�z��7�=�9&�:Y��?�I��V%LP��[�w7�U0Ĩ���M=�SX�x��{s A�|��=��1Y7ৌ�T��{Ǧ������4$�� x�]���.�Y���bb�W�J��@R%��.Y�����������~��T��F�����L�Y "U\��LV�n<�C�-s�f�}�x9l
���Ai9S��W5YM
t:G�1_�aqT��S��ED1;� �N�2yS�	�"�.�QAWj�������>I;Eܗ�h��a�л��L�Nm�:��*����r�[ǫ��}���Wz[��K�]��;� �𒑥J�e[�!*���D,�l�������t]dT�c��R�� -,��U�j_~4q�Jѩ	-)����F u��m��3w�cLF0	�y�	��MXmJ��{�4M!�p@�)H�Ü��t���%��q�+{*�e+����&�Cw��%�����r6Pf5��'�1|��Uw{S�A=SM��t�n��/i����*]�X�xnd�j����H^3�w	���-	j����ckv8F��4��UgU�l���O�1�4�ioIg��I/0�ї' �K��f��m	����Cػ���� �C�ι)�ހ
Gzj��F�8��d������r$��c?�y�9�Xܨ��#��}ȷ!64霔��o���.ѹ5ܴ{O'�4H{k�٦��3����uV�&�W�u��(y�V�TM��ŧWz���zj����X���r��w�*P�ae��&���2����@�a�fq	�� {���U�iCl�L+�_�uy)���Bk�����`4����]�(J�scp��c(�	���W� Y���-��'��B�7Ӻ̫�9����0�}�;W��\�Z�F�/��%*��3��M-�Y+��xT1'��n"?I��3�*������M8DL�-j��T(�`9�CtnE��
;�ߐI"w˘ݭB̽�/�Cof����B]�sw�e�$n��յ;��g����ؑ��t�\k�5(p��<_��k�~���)���:��<�|��./��:TSyʜ
�!����C�M5���a �Lm>N{�?�xdDe���)v2��`�<�_��bb8<k^6�w$`TJ�Fwd��$���[����>��;K�tV��MA�\��A�Zg@�3V������ -�՘/uq�����Q�� ����+r���X�W%���zP��]]t7Vv�D�m�w�Ӵ^���w!uAZ
5EgX^l�w����؀��բ�Ec�t�kJeЋ���Њ\
އy�ї?�U�0�q��y��6,6��+�p��-�&j[��K=C�) ���<b8���t'o��&W?˷���X���&ǁpP�7�8·0�?=��\��{.hl3��N4�y׸L��&,��"�;�8����#�I_�(�΂�q�s�2P��sN+m�ɧ�z��63��1� ����1��N�"@,~���E^���!����Kp���+!�;b=U�£^Q�^R@i��I��pqn��Y�P��B9~ =[����7R�)��)�[[7�7��$0h;��	�s�(e�ªQپլd'o16!�Y<+��n�I��֏l�e�Կb�|Fb_[v�N��VETBxG,�n3P�M*M�Y�����kۂ�]Po�.A��t���V+�8�#HjW�1�+hς�U��g<�Q	����f4
b�?��_�\C@�+2�a+G�{�9���c�0�)T�A�+z����X.�^�N�6ˠX���$h�A����8ωS���ͼ��o��z|�+<z��|W�CQ�2�4��C6��H�d��9sޘ�����}"��ͫ2 �1�c���4�J�.P��|"��D(5fv�&V��YU9�����98�'���(�^{�~�����o2��[�bԈ�:�o�����\/� _��)
B۰��`m�zم.8�@���1�/�S/-/�Տ8�+N�%�ʕٯe���?	j� ��"�ZuG��g��gl�/_]@�!	c� 7C��a#s���v��� D'bN���k3�b6�
��e��<�!7��^��q[	ɡ!��qa!%�����|9��q��[�\¸5	���4ᥠ��Kgu���ϼ�������u�Z|X�<e��/�.����@W19Y�@��Ħ��2��z���AR���y�#�Zs��Al�����,4��*Z���J}[q�6��"�Z�u>�`[8�F�L��R�t��^����#)'�_$[�v�k�O��E���g��E�wz��z?#g����>l�����	�����b"�3��O��zۉt�����j2���ٚS�R�{{W-��cQ219%`��e� ������=�V�o�D���2v��l5��X�#,��_e\O��-"m��IC��|�a�hP,�۰C*X�b����ٙ`M0ʅ'׭7�Н\;}�V����I�I��tFV�=/kex�MoW��ӳ��=�'�(�~{m3҄��FZ�)t,K�xSu�w�g����D��@/�����f�~* ��W=�Ρn���$�ȱ���7Ro�����"O@NR-�A���6yj�U���A�����LM����X�� D���N0�q�����	}+����l�0�����:�p��d��k���Lh���,@l`bg�@92UT<��l�-}:�1 ^:��S�4���(�14B�l��S��w1�ϒ�/�g��~+�u�~9�0߯NX pa ��ք:�gI�&���}_6����k���Z�\�!�@����ݭ�/d�?qDd1�J�����nEzA3��)jv?�2rL<梛���r:��<��\�X�u_����{3̣)�ュ�-
*�0V�{N�����97�b��φ.�^��s�������~&�D���>�Vx���Q�X�F�r��|�3����V�B�R���z���Ƈe�}��q(��b~;��(��fW��Cp?�W����C�����B��?�V����[�o���9y�o�u�m�g���Z}�ɐ���j��>A��Ļs��t��� ل^��|ڟz�=X����]"��|�9���2Q�c�IQ%E���C�"ۘs��ʎ�d�t���(F��5!=S�o�C��g���	
�vy::����Ѱ��X��[�RI��`BO�z�(�ïS�T�c�1˿�Dz�M��Ϻ��v�����h5�K�IVw_��|��s�O�1����bg9���5�@���63��z	���s�?�9
����#�q��)l;�N]g��V�2�k�
�,�f���)���^��k�m�Lc��̑���W�z��4���v#�x�ۭd�ȏU�f�4 �
��,X�sj�fȸ5*P0�Z�iF�	�q?��]��6d��_.��E��:O�ҵ��;Ng�k��tju��p������Y����z�W���z|�7-���)�L��R��z�����n���B����D��0��֤suo�{ت���Hy�8f7�9�FK�4����
�%�����z�Z��#��EM��K��
�Y�L�j���}X��j�@�t�Q��pm�L�"(P���o�t�4/bn���-iw������:�^�ze?�� ���ޅ�t�����6]��>��Q��Ras
�ء��y��"ƕ�g�6{�6�\i>v�@��aNM���K��P�Hb�kz VD^����ӗtZ� z�� ���V.)�)��r�pd���u����U][!�`�V��#�.8qz�b�����OC=4�.G�<�lk�.Yn�4D.z *p(�o�q\�#sŤ�[W-K�6��E�����
�Wq|WYWޫ������ݏ������ᕡ><���Mגx2+ @���,�ɰq���(��x��"��������}6�VF�˿�!xnz!Wqgj�"Y���kp
�����t ��3�uJ�1+��c�[�^NM:RN+Fa�WP���1�q��`[���ߏ��XӨ��Xs���z�S�aQ֖��li;�a�?��rD&ZЀ��U���_�����g��k��M{7!��ZD�ղ$��Y�J�pU!y�Jav�ڶc����\�~C�.���-��T�� ض*ZʡV)jXՈ����^��C�$$�m�=Aͫ��Ն��78s�_[�.dV���S�#nחE̲�JWx:�0-��z1�Ȯ
�Ȓ�'.��v@�R�ҁ�M���ά�-|7��,B�9�&jH	Z�y��|I��M���ե��g`�k,��N�k�Y�����(��a������d�ج��(<�	Q��.��hv�_MT��r�A5��P�X��z�%}ƔƐ�0Ė{�FX@�(�}:ua���������yv����A����^�Ѥ>�?t��r�h�����= �)���!]{Ls"n�|�lf',�A�&���-����s/'���z"+�#��������U��AP�zP%�P����^�̝�%��)8G��OA �T~������G�i�����`�\�&��:Q.Ȧ�X�$H�Y��'���Kf����*�m�{��Pׄ�fe�C�Z|`�����N���֨����e�l��W�E���$w�b1���F�H�:��\��@��]e�Tv���y�J'��P�=�%��������4G-Z[B�5�f�.��ҧ��4^y_���n�d��F�'d3��<�5�{	�;�h�[��bC	�������Id�t�|��+C�t�~p��r�����t/�_ya�Lg�K0�_�c�оxo��A�p���a��O�dܚ5n�޸�Z'g�i��{cWf�tr��ɔ��7D�1�$1��=�2C��a-]h)���hL}��Y�g'a�1��㎏��/n�9�����#
�N�L[^Ro�9�0
�F�9+�BFv4- !-f,�\U��/ɘ�K�i�����HH�+B�j�I_@�����>����UV��%�N��MEz�[YZZ��uQ��������
�R�h�~c��t��>Y���3U��ҫ6���:ؽ7xc�\��v@��Ui�� ݂J�q��2D�(y��<�نz�ɂ��qR��]"v���.���;����Lf��43@��M������RA�kݒw�lV^�+��*�寳�ϼ�k����A+Ob���%TG>G�
&m!���As�j��6���sJ��L8{<Ѫ�l����~=:(�S�T���s{)�]*�*�=�S��?�!z�Fz��H�6X�s�&r�e�cz~�d݄�p�w�f+��x���[�oO������j��a9zæ�Z l��g�(� �,�%U\r��0���<��{�5_�im:ka���2�3�S!���gY�G+Hz	��=�K�xN����~�}`i��r;����)�.�yL���`+�F9-?C��R���zt�4��� ���ؘ���^A01�;)[9=�F ��g�Iԅ"��A|�D��L<������]�i�IY����r3���]Nj���b�P�)J]0~���Q�Mq�j:帱���`�"�s��Tב�gT�t���4q������>�ǞZ34^��H��Ze&�.����s��2c��y(�V�A���ƚ��u����6��������0�C�܃��5��e8�P��7���f���%�#���� (��-�4�����o鏸~�S8��\h�R�Z�`�|�>���o�G�ֺ�K�$�b�Q�%^��=D]0�G��m�2��G�w�؊qO|%]��LW���j����H�B�ϨB��ި{(XUPZDN�8^Z��e�֡���/��3f0�!�х�5��8��1�_���/����e>��- <=B�}:�eᔥ��H*����,��=5m�ov���xjF�ҡj&�����=�O���3��;%5A��W�1F'�����m�f0`��"M~���t]�=r�&��OVш~�����Z�g����˥@ -�p��ӤP�cq�$�����U:@'/���l#e8�|U1���`�G=ꊍ3l�4H�-�0��g�RgPs�P���L��PG���0���S3q�r��⍛]����"�7<Z���x����I�����1���"x{��*#M��:���rq)�v�H����`��r��M���7j_�B�*�q�TO}b�mzu"��P��+�Ai�F��tMԏP���ظf
��V���O:�湺�<7�����h���q����8c�
w��uNu�Fqa	V��o�/k�"׉
C#�!f��wT�{��P�t7?z2��Z<���*��㳀���¬{~��7ZCׂE�XU�%&$�#݇zv��z�h�AG�5!i��$_�J���>�W{�%+�F�R�<|u:�`����fҝ�yMD�iۿ�AE�K<��<����.}�C��!��]����O�����D*�?J�.l�����%5Z"�,$�PIn��g�xbR�,�i �
C���d��cTg�4��9]��C+���0k� 4�rl�Sd�D�{�����f!ߡ�R�0O҉R���\��sB�"�ǣ���M���uGT֔�d�T��R���)L�+{�,��W��p����,�q�.�?�R^3W.�D�wWa:��{�vz�7⛫i�6\ֵH���^R�rD��^h�|��*��9$;-�;�>�0��58ʾWN�W���, u��]�EG�ѹ�d�g-{H��w��	ͅ�Jhޤ L.n�Ѓ����H�r��Xz�UH��PR�c۸Hg������&p�e呋G<��]��C��g�iSZ��h��^H1�!��p�=��S�_��>��E�D_7
����Cp����y�$�e}���^6!9XwQ>.&Ӂ���ꦨ��/[#�
�﶐�A��P�fϹ�a���0ƛ͛��9?�Oky��h8������熖����f�"���ۈ8�;z�Vˮ��\����X�5,^�k�Y;���>�b�欀�J���}mm��������&M���=W�>J��<z!:���Z�ROL؉ErG����^�+Y<�F��H0kR�L������vǇ��
��YS�h���N>�D��`�eB߱ ~K�A/������Y.+�g��!t�#%M������SS�I�z�-&��j���n)M�ɻ��(I�w��&�K�|��g*3�5�VQq�PM�ԉX�t�xF�0�6��11�����Y��k���J��p�U!���q���cp��ګ�oJ:��X��*��,�d>e�I��;$�)Gs)�1�0!҄t�' �U���̤ZF9���If�J��B���1��NA@�0u���Ķf3w�p����1��0+E$(�h���-A���U�b�$��&�fR��G$%���ԝC���UK�����$-\�	�-򥛳;J�%NI`�ͼ
>�F-^���L����L)��(5��C��?���Z6"����J�w--�Z�p�������5����I�b���(�[ޕv3+��F\;6wޘ�*J��,�e�{?���%���&����5�Y��((��W��a'%���ɝ�I�����J�lc�ѵm��	[.�Y9q��6�M��hI�N�Łr����AC����|�����k��������Gt������8�P1^��D����@����}�=+k���,Z\I�t閂�����	k7x$s�Cz��&����)�[��6誗WL�������_��)L�OU|5�Y������fr�fFT��(�
�Gw��__��qܖ����v�/@V��P�])^H���{�B�0��}�"x���D��:���i4�o�]�i��ۨ������Ǜ�M
�B0�a	t�x"(�?ΰ�]�ͫ O�D;&ãXr4g*��>S���!uUt}wPGq4 X��KS�r�����t-�V���O�D������ȃKf�6���h�5���b��?�7w�����]F���(��:��LF��Rn�=.��Z�VLz�I�%d��]�q��gi5�K�����ν�m.h-�.��FA��� ��'V��K�@v
'����q�)�ۗy�4�q�����o@�}��/��'j)����Ha�L��V�GL���Z��1��wu����c���,&��>��d�V�w��
��"H,�ؙ�n��TZP�@>j��S�[γ����j�X�~|?�uV"r�y���X�h�x�0�+�^Ɯ�տ1��S�Z���ы\B����,B^śj���٩�ړ��!�'�W����<y�"�~�N�@ƼN��7µ�
�S�Z��㹃����vwh,�-B��Z�9��-�牂?+A�����yR�4���C�([����� =�E���R@�B�I�L�o/WލF����?�T���0]O;��A���7U�Z�MX�$5b{y�ҭ"x8�ԇւ�_a`a�Hc0�&@�U�AS
����Y�#�����j�������`
��	Xc,�m븉�۫+�(j�D�љ�)_D}��(-��El��Ae����P�&vj����!�k��/k�q@~&�;�7ü1|�!fv.y<�V��1��u.��f�t����V�Tr��&F-�mP�L���-���~ d�G
 j�t7�D�7��4\�v�f|x5)��	uc��9c�}�@Uxe��>R���t��B�TƐ!�/o M���^(��I]��Y���jj�f�$�k~􂤫���[�3�d�@�]��k���28����i!���&lK�Pg|��9�ĵo-u:r�$PD�VT�Z��N�S��'�x�FcGrL~��e��s�")ԫSC�΄y�<4���<J�%���a,�R}pQ-yc؇ .ؼ�N�e�/���_VS+��3\�0�ö2[���vt$���J�������+�0G)�cE�&X��ڈ}M�]xs��k��o# ����Z�]�^��z$YBv�uHg�5ns�W=�������eE~O� �G�+�v��
��|��<���Z��QnQ�.ŝ����ЯEB�
Hc����]bq�	 +��F[4B�~��}�,Ǹ+?Ш���c�o���n���:�jG���ʄ}JC�/d��i�_O���)�S�U].K�ϯ��dQn�`S/�ou L�;�w]��3u73l���p�NS�ه`6#i�*g(��>�_Sȓ��|Oh�*�F� �Їl���'���	�1��/���bҸ����"V��~|W3T��Ay	 �%��w1�㳔����{Gr�/2k��v�xx�n�?�i6Y�]��Pk�V+2�O���~f��	R.�D��,"��3����(�����4y�hCR�%��d��%���ǎxb �^�O>=����s��?R�o��΄��b��D�������ߵ��A�-�𜖪H��+ �K�4?�RW���25R ź�_S`̈́d���,��@�����0 ym��� ���OѪ�[�Q)) �v�i����oք�Y-&*F��+��Y)��A����8��� 뙿�s�X]t��T��y'�؅��m=2g��C��p��L]n�'S�n�z �ޫ���^h����e�����2s�>�n0B�SE�d1���_�F�7%.�|�M���R�W��<r�S�PH<������.�ĥ�9Ŀ҉U�K3Vh읹��O/W�����Q�����y����uDM(�%~���
JM1*�Gս� ���.��?ҷ� y f��'�˨����uo���n١���=�%¹i;
��� N� �;��N��0K^�[<����A��rB�oT#	_������qF���BBih�&���+�f���p8����������Q;�|gI�_���¥��S #D�jY�Le��ά��}�n��~Xi@�τ��c�l�BRtm�|�^(���|Ę����6�j��:�9���mz��p�w!�է�����������jB�S�!>��D����}�� ��S��`�U���ϝsn��w�VyK�����黗p!��Ç�?a]ʟ�.C?hGg��~��h�e�� ��g1�(�i�[�s��L�$˃&m���Y;G�d�<z�;��|��_�y�h(��-���s`���gvQ��}����m4���困*���"�Lq��+P��?�GXm��`��`�Q�{��.�yְ���ٓ$'B66.R�&��1X<dQey�\W�TUO��/�e �)|�9�^W�t��)f)XlQ�}�����"�i9,$cN\&E�i�a��BQy�6h�������Q*!]{�jp�9�8JKY�K�c��.�������s�)�M��3��e^������vS�+A�Q�7E�Er���d���4��;�'^�׾*P���"[,O�� �'�����I�S�U%X��f�.����9��~��(ܐ�W�e�5�8����m�3scN�i��~Jr�Ϙ#*����,1���[��LE�ѝ�(;�ң#WRf�l闬�J*�	��N�[�����eL�'o��G �m���������ߍ����8�c�W�][80��ʄ��Q�-��׏��!�@Wy{�����Ӫ�bkc�s���� �T��3���Ѐ���͑�AȆb6<���U�Ѓ�F^��:nׁ:�[#��M:u�$`+v��1������̀9��^��Q����FGӀ�Ө
�~�<���&<�@i�)~�hL�Jl3	Вv#���>�D�^�J���M��-H$|���H7�<\��&:a=����]����/�/����W3Y�K(�i)A����eo�q :_Gp{�j�tf��#����Q�p��Xs���6�ʀ�?���]ѽ��c��]�
%��D�rd��8e]��.�"�҅�&��H~q�}���A��M�p����<ߊ�'�6��*9���9��9M����'9g�R��nz'��t3�|@�P��o�������jx��3
�2xߓ2��m��e�i`f�U.����M@�BuGd\�������4X�hg�-�9m>�<�g�Et��-��a_��<��7(G��;�ő;����8:�'���j��zD���w��EȌ����x� #���M��{�\K5��9.�1���n���VG�FI��3�^����k�n2+r6y#����<�b_�"Q�(������\Ff!�*T�YjJ<��h8�}.�lqpQ[�\���+�!��Z�t��MA�I��O�1ӛ%y�!��y�R��>���eh�4`�(%�Z�:z��I��c�*��h(�ށ�2���Q� �ܼ����b��l'}��9������e��T{�2����́�X�%j�������6!��pg=� ��Ξ�xzs���Cj�E�JS5�̃���)��[�N��@�
dpԄ������	,��t�S�]����w��� e`+8����l�ӏ�]f�B�?�0f"a+��&�ع��z;�i�;�|S�l��n\f��~�������m����*�ea���!�̻��%�T����VٻR�d�}6<�L�w�7�"c�z'��� ��IrJv������J`�2t�OZ�)�գp��j�҆�IH�Ur�D�D��F+�X견J�䣢q�_|n+9�&��뵪��=���v�Ssb�[(\��++��>^A�^�H��n�7�!��mIL�!�����O�(��!ĠI�LS�W�S��m�K\�a z\��jk�����rβS_��c
F(�q��t�w�:���8����ĺ7B���ă|7��mk�@lC�������ޱ�� ����h-f(����
�gm�_��f�ZfΗ��G��RPzR�↛������b	e��
gc����茠 >��ۺ���� bS�i�8��'�&qE��gK��K�W�B���Į��Ġ�fݠ����>'�g�`>���Q��wr���Oo�յy6A�3j��扙���	Rʙo��TؤWW%�r�߮������8�m�
�ۈ#���q�R�K{C�Z��|T����'ƌZ�_�cܬ,$�n]=�L����>r�s>b�Y8	���������n$5�����;!j�����i;aQH�^pS'N¬��s83��f��� �n�ke(�	n��^#b���K�u��G2JWX�jc�r�,J7�g%K��9�Oh�-0���aTL
�ʓ����[��ģ��y�LDv�����Ƃ����94g6>�}�5��Q���O�vr��s#�l����=!n��p�*)6�)=��>��t.�m�k=tB�K#Bn���eͺ2�戜�I9裥�f� "�+������ �8[�JZ"�����;���I��v��W�TgV,����b����Y�(�c_���D�rܤ;;z�o��4Hm"yKFn�I�!��z��|A�O��O��dў�'�����V51|�&�c�OT��I�d?���G�n��MPPc�#KFK�*V�MM?�sQ􈤹�t�Z�-���n�6�2�����_��1�K�:=�GG�7�Ȉ-(u��ڲiD̀��((�n̺&�)_�H�ˁv��]����0ۊ�J�X��c���X"'YS���� 蹢���$��^o3���>@3�}�c�O�o�)�yIQ��i�RR�yY�h�4G	ԙ�����J��CX��5�Dlr�X��'�	��I��X$D�6��sN�Kþ3�"��+;�W��p)E����ѻB��Y{���ţ�GM,i��'�i�lUʮ�u���W�,#�0s�ٴ)L!�G�|ɡ�	��O��l>{)c�<rg
 �EТ�zY�x�{2�&�X���+
*�w�e	��'���0��r��25R���|�9�Z\�g�Ur>&
�:�2�پa�~�����&:���T`u��A����W����1v�N�;��ȋ������� YԼ�<���[�ĵMEwvU�#��j^J����i�C�� �V2��HP\*����+!)���+�V�J<T�!=ߎ�uc
v�k�|��W��JZ�S�Ƨ��=Ƕ��^�A����빧b�e�5cd�T�pc�[m7��G
	�ԄN�<����ݯ�_��ݡh_����𢦣���OT'��,����i���^��>�.t�9l�C�=^�Loq����岾����&�.XR�3�&@������rV�$�^��y �\�h�	����K�Ɠ�K_�J����Z��k[-�u ��ZA�G��F��,���~ �v�h�����n�K��ĕO�h��!^�����B0����p�`N��u��XS��_�$��<[�����]yW������?�۠!W"�����]^���A[s4:��r-�c�Vj�.�� 3�y��%�:��C_E��_E��(Uu^T6C���r�@��IIJ�$�%5���KQ ��`|���3~�Z|�eN0�?a����!#��,�� �h�LR.����W�W������wJ�lҢ���g@��O-ĥ!���=���SKχ�r� ,BB6�#���ᐜٟ��Sl�gy�	ʹSݔx�L��t���y�l�n�Q;��G����pE�O|��j#!w��ya���X�b\��f�s�)Qy�Ɂ�T��х�0������|�=8K0�#�hKӎ͓M���hd�U�a&2;J�%y�#a�+¬0�T�_��؋z�ݰY�y��lIG� ���5���׼��g�}�Z���8cÖ#W1�=xVf�lK�U���
j wWװ�)�8��Eb�w� �G��=qQ?q?J�k]���fBCD�+u�#]؋i� 2�]�j�%�T�j!쥲�`K@�����"g�aTSX��R䗐^�e��.���(X�,jc�eWx���7QN�Og�xh�.[h�G0ȸ�8uBo��~�Z,&W�H�[B"��u�".�5v}%��K7�⍨��tш4�P�A���!��C���Ă��C�G�\`g����1��u��,ס�&A
�,`J��uo�Knl�xe�q+�agt,Ǻ�v���[{;wEA�ۘ�C��A`?h�!�$��;�j�F�pOgը�,c���c��
)���$�i.�O�BQ�<�絎H`�#db{����3����o����6�
��A��A�����Ƃl�0�S�47�k�I��Dø0�XxGǚk�f�������zR�B�d��L�7�gQ^G�0�cw�-����1bٝg<�fqa#��'�:��[}�c���wѵ!���Z:`<[@e��T���(��W��BA௬'_'1���LB��S�U�p�l��ܭ ������&�`F(���e9h����/��f1��B���x��,��c8Z]�� �xE�n�G0x��#�F�Y��5ܦ�#r1� ՈN�yΆ}_�� /��"-�sh	����O�W��ǡQ<��ޡ L�L ��	Y1�����m��]T�z�m�ؐ��@n0�������w�B��y[����&�,!\3�kGau�����'=9d�����s��,s��}tՆ:D����i�P�����њa�u)w�����
�����`�S1p��qD}*��#0�Bլ�7/�����a"s�!qa�v��O�v�OR�;�y��X��Cy�f�����ȠV��bs�1/��i�]�G"U�Ȅ�	ͼ�������pX׺�����)�~�Ӫrpb/B�EWK������$�2�$�_�Sj}F�bEܔ	�|{�Rw��o.k������U������뢚tUH�cB雓D���Ne�y����"f�.0�Ŋ����G� �U%;�־��=GFoN��S������M�\u3�Kn£��~���~W��ϟ'�b�Nj���0�8\=J�R)HW�)'�T�&<��pzB�{.� qi}���s�W��X�������e��P�O𫏩L
�"�mx0�-�`���-Y `��b��~��M��\|�O#j~'���*��]��&B	��BC�f�H�$�-���niG�� (��Vv�q�s�M�T/����vN.���|�䎓z�9�f��Vb���e��)�أ�BFǨc�X@ȿ��i~�t��Ę�4��B��m]3��>��ϖ�>�qi�����r�y�b�E3&f�d�Y��T'} gx �~I�k3X���qm�f*��j@�/s
����6��L2����>�Jк;#1��Q��)ꅧ��[��oE�Uxg?�	s��$q�x��` ڊ<����n�Ŭ㩆&e���y<VU��H�KW�^%�C1�^�P�ak�;Q���aV>�d��Hڽl�C����a�H%�J�{�k�T�*5y�Q�O�{�ta!��4�<%?ZZga&�h3��!bq�!)->�sW%8���ރ�+3����F�f.���	��ᧈ�����ٌ!2�ua�?H+�� Mժ:��|�O,6Қ�~��@i����XnR����z+���3�S���y��CJ���Q*NU0#rU����rX�y�4֬^K�x�a]ŏn�:��!'
@�~�@����y	�՟�$�V�N���K%&l��E3Y�Q��>��y);Y<�3�9�XEh^Iz:�8z��B��-M���q�n�%�p��M��>CT8β�-��+!�}�5|�&�F�E��c#ϴ����&��doH�V�� Z`�� �Uv$m�S�Y|�}Cw�6�L r�C�a�%sq�V�:W�E�!을ʹ���vxS��΢����٭[k�Hf�Ŭ=/��FA:�i�b��Q���HG8d�F8�'"�eBd�姴9�7ԱN'*��s̏�˛���H�`(6-�I}���I�mz�ՙ�f���^9��'�(��Do�~���*Mr<�Bҝ�>�j������EL`!Ǐ)�w��5w7��\�&�'Io���}_�}���eS��"�"��v�g����af�b�饚��C^C"������^;��_^s��k�iYXÌ[���Ql����N$t��P����������*���:@
��:�h��VŘ}���_$�4-?%�X�"�ǈC�*�ԇ�p�qKlq�UIE�#�<�e�r�����f�%��垔���Pmz)�ԏl�k����w�������
� ���Bq�(��#y��Z>TL��YU^߫m�ɀ�5ԝ�=\�1q�	�D��V�y�i*��I�3�vx�o�-w�vu��J��;�]��X;E m�ˡ��P��O�"`����{ӳLK���\]������R��J��ߕ9hc�z�}^�j�����z��݌"���V_!�D��c�(:Y��t��L^}���P�9��WG3d1�.|�Cn6�y��]|R?�ae.�(��q���X)qt�1�6�
Y���c��	�7��Ѳޕ 2B�,�USJMI� �s8fZ���#�0�'՞+�|<���vq�B@Y#v�ҟB<���q��u�2���l�t����8R'�(���J���(3,�4�V
�����ն�$b$4�����7�Z���B-o��ܒk�w�@Z4�� ��G6bR�P����.l��Ի7I�3��#��	a�^C�Q�%��Z"����F荸#�@&�V�h�?Uj"��-3��A|�0+��[�Ǎ�]<��u�Ƥi��3L|��O�K��;4ѴǼ@�Y�c;���]��!8&��K8��]EW��T�Z=Π������۰5g^"�a�0_��c�-���_��G���j��6���j�L��H�����z��+�ɷ]ӳ��+m��%}]ԋ�f�=�c�_�3����9��b�XvE�a�lUUD��:�&�|hA{n �".��=�}�%P���U�M����ÿ�A e�x���,���$���j�@M�N��^�#~�R�F�/��բ����;�_Wp9t���~�:���a����S	Z/w���]��Â�}�8�{�Gx��}{DWF!�2�r��w��*�D8t��g����Q�k������s��'c�,O� Rp�~;���7�':����+c^�l���ʏ[!?���FJ�p�@�����־2�\G?`�)�[��N�/y�wW�&���)�c@������ ���#AL�Bd�Pv�ni���������\"K�2;�=ݽ�j�,~ଶ_t'W��:��&��mH�A�#e�=_�K�n?ha�9Q�G�W��k!�
k�:ž={���c��H�����Z����2���2_�gWU��竗��)['-omJ`��G�Ozk|����k�����Z��53i��^^*ݏ��Q�����:[R���r���W��w�i޷��a�5�ʄ���T�[R�Õ���F����7��������yS��g��DdJ�F����:b�HH|t��MШ��X�с�dr^@^�V�J~T�oFT�V@%�(:bG-*���V�>g�7�T- �Y*��Dl�*�h���!N��KqŖ1�J�Z�(}�ބ�w�H��xT���%R�i�SH*V.�Tܽљ�D#�dߖx+rxfyYG���f��f��q�M�������C=������*�[����]n&�J��n�����_}Xԍ�\�o��l��igQ!�̀A{�BM��B3l��=��q���3Z���)�%Օ�����&>x>ŭ����$x��Ĕ�l��p[�L��5"u:zض�N6�V�0I�Y�����SU6|<:�P���e�z�^�]���H��+~p�g�04�)fp�k+䖡D�̆�Z���p��B�P�~"�W"�i�V�K����������f���<����!��3W�R��L���p�y�/�6��c���M�^��a��*E���:W�}��"S�"[}>'
��P�+��n;&���)g�����PY�Y8����zP=�w{�)�-�oA���w�q��<�)b� '�(<	8��!\q�`����x�<�$����~�n��:�"*,q�](	��r���~�8�gL.�	(���8�EQ>&)uçfm��Ee��`WP����`e����xDo?R_a�'� $'m��4/�p��9a��a��I�|z�d��G����u��