-----------------------------------------------------------------------------
--
--    COMMERCIAL IN CONFIDENCE
--    Copyright (c) Commsonic Ltd, 2010
--
--    Commsonic Ltd,
--    St. Johns Innovation Park, Cowley Road, Cambridge, CB4 0WS, England
--
--    E-mail    : info@commsonic.com
--    Telephone : +44 (0) 1223 421845
--
--
--    Project name          : ARCHIE, v@project.version@ (@project.revision@)
--    Product ID code(s)    : CMS0041, CMS0042
--    Block description     : DVB-T2 Modulator.
--
-----------------------------------------------------------------------------


 
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_arith.ALL;


PACKAGE BODY cms0041_config IS
  PROCEDURE user_cms0041_config(VARIABLE v_config : INOUT r_cms0041_config) IS BEGIN
  END user_cms0041_config;
END cms0041_config;

 
 
