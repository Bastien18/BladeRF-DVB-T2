// nios_system.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module nios_system (
		output wire        ad9361_adc_i0_enable,            //        ad9361_adc_i0.enable
		output wire        ad9361_adc_i0_valid,             //                     .valid
		output wire [15:0] ad9361_adc_i0_data,              //                     .data
		output wire        ad9361_adc_i1_enable,            //        ad9361_adc_i1.enable
		output wire        ad9361_adc_i1_valid,             //                     .valid
		output wire [15:0] ad9361_adc_i1_data,              //                     .data
		input  wire        ad9361_adc_overflow_ovf,         //  ad9361_adc_overflow.ovf
		output wire        ad9361_adc_q0_enable,            //        ad9361_adc_q0.enable
		output wire        ad9361_adc_q0_valid,             //                     .valid
		output wire [15:0] ad9361_adc_q0_data,              //                     .data
		output wire        ad9361_adc_q1_enable,            //        ad9361_adc_q1.enable
		output wire        ad9361_adc_q1_valid,             //                     .valid
		output wire [15:0] ad9361_adc_q1_data,              //                     .data
		input  wire        ad9361_adc_underflow_unf,        // ad9361_adc_underflow.unf
		output wire        ad9361_dac_i0_enable,            //        ad9361_dac_i0.enable
		output wire        ad9361_dac_i0_valid,             //                     .valid
		input  wire [15:0] ad9361_dac_i0_data,              //                     .data
		output wire        ad9361_dac_i1_enable,            //        ad9361_dac_i1.enable
		output wire        ad9361_dac_i1_valid,             //                     .valid
		input  wire [15:0] ad9361_dac_i1_data,              //                     .data
		input  wire        ad9361_dac_overflow_ovf,         //  ad9361_dac_overflow.ovf
		output wire        ad9361_dac_q0_enable,            //        ad9361_dac_q0.enable
		output wire        ad9361_dac_q0_valid,             //                     .valid
		input  wire [15:0] ad9361_dac_q0_data,              //                     .data
		output wire        ad9361_dac_q1_enable,            //        ad9361_dac_q1.enable
		output wire        ad9361_dac_q1_valid,             //                     .valid
		input  wire [15:0] ad9361_dac_q1_data,              //                     .data
		input  wire        ad9361_dac_sync_in_sync,         //   ad9361_dac_sync_in.sync
		output wire        ad9361_dac_sync_out_sync,        //  ad9361_dac_sync_out.sync
		input  wire        ad9361_dac_underflow_unf,        // ad9361_dac_underflow.unf
		output wire        ad9361_data_clock_clk,           //    ad9361_data_clock.clk
		output wire        ad9361_data_reset_reset,         //    ad9361_data_reset.reset
		input  wire        ad9361_device_if_rx_clk_in_p,    //     ad9361_device_if.rx_clk_in_p
		input  wire        ad9361_device_if_rx_clk_in_n,    //                     .rx_clk_in_n
		input  wire        ad9361_device_if_rx_frame_in_p,  //                     .rx_frame_in_p
		input  wire        ad9361_device_if_rx_frame_in_n,  //                     .rx_frame_in_n
		input  wire [5:0]  ad9361_device_if_rx_data_in_p,   //                     .rx_data_in_p
		input  wire [5:0]  ad9361_device_if_rx_data_in_n,   //                     .rx_data_in_n
		output wire        ad9361_device_if_tx_clk_out_p,   //                     .tx_clk_out_p
		output wire        ad9361_device_if_tx_clk_out_n,   //                     .tx_clk_out_n
		output wire        ad9361_device_if_tx_frame_out_p, //                     .tx_frame_out_p
		output wire        ad9361_device_if_tx_frame_out_n, //                     .tx_frame_out_n
		output wire [5:0]  ad9361_device_if_tx_data_out_p,  //                     .tx_data_out_p
		output wire [5:0]  ad9361_device_if_tx_data_out_n,  //                     .tx_data_out_n
		input  wire [1:0]  arbiter_request,                 //              arbiter.request
		output wire [1:0]  arbiter_granted,                 //                     .granted
		input  wire [1:0]  arbiter_ack,                     //                     .ack
		input  wire        clk_clk,                         //                  clk.clk
		input  wire        command_serial_in,               //              command.serial_in
		output wire        command_serial_out,              //                     .serial_out
		input  wire        dac_MISO,                        //                  dac.MISO
		output wire        dac_MOSI,                        //                     .MOSI
		output wire        dac_SCLK,                        //                     .SCLK
		output wire [1:0]  dac_SS_n,                        //                     .SS_n
		input  wire [31:0] gpio_in_port,                    //                 gpio.in_port
		output wire [31:0] gpio_out_port,                   //                     .out_port
		input  wire [31:0] gpio_rffe_0_in_port,             //          gpio_rffe_0.in_port
		output wire [31:0] gpio_rffe_0_out_port,            //                     .out_port
		output wire        oc_i2c_scl_pad_o,                //               oc_i2c.scl_pad_o
		output wire        oc_i2c_scl_padoen_o,             //                     .scl_padoen_o
		input  wire        oc_i2c_sda_pad_i,                //                     .sda_pad_i
		output wire        oc_i2c_sda_pad_o,                //                     .sda_pad_o
		output wire        oc_i2c_sda_padoen_o,             //                     .sda_padoen_o
		input  wire        oc_i2c_arst_i,                   //                     .arst_i
		input  wire        oc_i2c_scl_pad_i,                //                     .scl_pad_i
		input  wire        reset_reset_n,                   //                reset.reset_n
		input  wire        rx_tamer_ts_sync_in,             //             rx_tamer.ts_sync_in
		output wire        rx_tamer_ts_sync_out,            //                     .ts_sync_out
		input  wire        rx_tamer_ts_pps,                 //                     .ts_pps
		input  wire        rx_tamer_ts_clock,               //                     .ts_clock
		input  wire        rx_tamer_ts_reset,               //                     .ts_reset
		output wire [63:0] rx_tamer_ts_time,                //                     .ts_time
		input  wire [7:0]  rx_trigger_ctl_in_port,          //       rx_trigger_ctl.in_port
		output wire [7:0]  rx_trigger_ctl_out_port,         //                     .out_port
		input  wire        spi_MISO,                        //                  spi.MISO
		output wire        spi_MOSI,                        //                     .MOSI
		output wire        spi_SCLK,                        //                     .SCLK
		output wire        spi_SS_n,                        //                     .SS_n
		input  wire        tx_tamer_ts_sync_in,             //             tx_tamer.ts_sync_in
		output wire        tx_tamer_ts_sync_out,            //                     .ts_sync_out
		input  wire        tx_tamer_ts_pps,                 //                     .ts_pps
		input  wire        tx_tamer_ts_clock,               //                     .ts_clock
		input  wire        tx_tamer_ts_reset,               //                     .ts_reset
		output wire [63:0] tx_tamer_ts_time,                //                     .ts_time
		input  wire [7:0]  tx_trigger_ctl_in_port,          //       tx_trigger_ctl.in_port
		output wire [7:0]  tx_trigger_ctl_out_port,         //                     .out_port
		input  wire        wbm_wb_clk_i,                    //                  wbm.wb_clk_i
		input  wire        wbm_wb_rst_i,                    //                     .wb_rst_i
		output wire [31:0] wbm_wb_adr_o,                    //                     .wb_adr_o
		output wire [31:0] wbm_wb_dat_o,                    //                     .wb_dat_o
		input  wire [31:0] wbm_wb_dat_i,                    //                     .wb_dat_i
		output wire        wbm_wb_we_o,                     //                     .wb_we_o
		output wire        wbm_wb_sel_o,                    //                     .wb_sel_o
		output wire        wbm_wb_stb_o,                    //                     .wb_stb_o
		input  wire        wbm_wb_ack_i,                    //                     .wb_ack_i
		output wire        wbm_wb_cyc_o,                    //                     .wb_cyc_o
		input  wire [31:0] xb_gpio_in_port,                 //              xb_gpio.in_port
		output wire [31:0] xb_gpio_out_port,                //                     .out_port
		output wire [31:0] xb_gpio_dir_export               //          xb_gpio_dir.export
	);

	wire  [31:0] nios2_data_master_readdata;                                        // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                     // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                     // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [28:0] nios2_data_master_address;                                         // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                      // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                            // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                           // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                       // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                 // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                              // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [17:0] nios2_instruction_master_address;                                  // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                     // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_command_uart_avalon_slave_readdata;              // command_uart:dout -> mm_interconnect_0:command_uart_avalon_slave_readdata
	wire         mm_interconnect_0_command_uart_avalon_slave_waitrequest;           // command_uart:waitreq -> mm_interconnect_0:command_uart_avalon_slave_waitrequest
	wire   [4:0] mm_interconnect_0_command_uart_avalon_slave_address;               // mm_interconnect_0:command_uart_avalon_slave_address -> command_uart:addr
	wire         mm_interconnect_0_command_uart_avalon_slave_read;                  // mm_interconnect_0:command_uart_avalon_slave_read -> command_uart:read
	wire         mm_interconnect_0_command_uart_avalon_slave_readdatavalid;         // command_uart:readack -> mm_interconnect_0:command_uart_avalon_slave_readdatavalid
	wire         mm_interconnect_0_command_uart_avalon_slave_write;                 // mm_interconnect_0:command_uart_avalon_slave_write -> command_uart:write
	wire  [31:0] mm_interconnect_0_command_uart_avalon_slave_writedata;             // mm_interconnect_0:command_uart_avalon_slave_writedata -> command_uart:din
	wire   [7:0] mm_interconnect_0_rx_tamer_avalon_slave_0_readdata;                // rx_tamer:dout -> mm_interconnect_0:rx_tamer_avalon_slave_0_readdata
	wire         mm_interconnect_0_rx_tamer_avalon_slave_0_waitrequest;             // rx_tamer:waitreq -> mm_interconnect_0:rx_tamer_avalon_slave_0_waitrequest
	wire   [4:0] mm_interconnect_0_rx_tamer_avalon_slave_0_address;                 // mm_interconnect_0:rx_tamer_avalon_slave_0_address -> rx_tamer:addr
	wire         mm_interconnect_0_rx_tamer_avalon_slave_0_read;                    // mm_interconnect_0:rx_tamer_avalon_slave_0_read -> rx_tamer:read
	wire         mm_interconnect_0_rx_tamer_avalon_slave_0_readdatavalid;           // rx_tamer:readack -> mm_interconnect_0:rx_tamer_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_tamer_avalon_slave_0_write;                   // mm_interconnect_0:rx_tamer_avalon_slave_0_write -> rx_tamer:write
	wire   [7:0] mm_interconnect_0_rx_tamer_avalon_slave_0_writedata;               // mm_interconnect_0:rx_tamer_avalon_slave_0_writedata -> rx_tamer:din
	wire   [7:0] mm_interconnect_0_tx_tamer_avalon_slave_0_readdata;                // tx_tamer:dout -> mm_interconnect_0:tx_tamer_avalon_slave_0_readdata
	wire         mm_interconnect_0_tx_tamer_avalon_slave_0_waitrequest;             // tx_tamer:waitreq -> mm_interconnect_0:tx_tamer_avalon_slave_0_waitrequest
	wire   [4:0] mm_interconnect_0_tx_tamer_avalon_slave_0_address;                 // mm_interconnect_0:tx_tamer_avalon_slave_0_address -> tx_tamer:addr
	wire         mm_interconnect_0_tx_tamer_avalon_slave_0_read;                    // mm_interconnect_0:tx_tamer_avalon_slave_0_read -> tx_tamer:read
	wire         mm_interconnect_0_tx_tamer_avalon_slave_0_readdatavalid;           // tx_tamer:readack -> mm_interconnect_0:tx_tamer_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_tamer_avalon_slave_0_write;                   // mm_interconnect_0:tx_tamer_avalon_slave_0_write -> tx_tamer:write
	wire   [7:0] mm_interconnect_0_tx_tamer_avalon_slave_0_writedata;               // mm_interconnect_0:tx_tamer_avalon_slave_0_writedata -> tx_tamer:din
	wire  [31:0] mm_interconnect_0_wishbone_master_0_avalon_slave_0_readdata;       // wishbone_master_0:dout -> mm_interconnect_0:wishbone_master_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_wishbone_master_0_avalon_slave_0_waitrequest;    // wishbone_master_0:waitreq -> mm_interconnect_0:wishbone_master_0_avalon_slave_0_waitrequest
	wire  [23:0] mm_interconnect_0_wishbone_master_0_avalon_slave_0_address;        // mm_interconnect_0:wishbone_master_0_avalon_slave_0_address -> wishbone_master_0:addr
	wire         mm_interconnect_0_wishbone_master_0_avalon_slave_0_read;           // mm_interconnect_0:wishbone_master_0_avalon_slave_0_read -> wishbone_master_0:read
	wire         mm_interconnect_0_wishbone_master_0_avalon_slave_0_readdatavalid;  // wishbone_master_0:readack -> mm_interconnect_0:wishbone_master_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_wishbone_master_0_avalon_slave_0_write;          // mm_interconnect_0:wishbone_master_0_avalon_slave_0_write -> wishbone_master_0:write
	wire  [31:0] mm_interconnect_0_wishbone_master_0_avalon_slave_0_writedata;      // mm_interconnect_0:wishbone_master_0_avalon_slave_0_writedata -> wishbone_master_0:din
	wire   [7:0] mm_interconnect_0_arbiter_0_avalon_slave_0_readdata;               // arbiter_0:dout -> mm_interconnect_0:arbiter_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_arbiter_0_avalon_slave_0_waitrequest;            // arbiter_0:waitreq -> mm_interconnect_0:arbiter_0_avalon_slave_0_waitrequest
	wire   [4:0] mm_interconnect_0_arbiter_0_avalon_slave_0_address;                // mm_interconnect_0:arbiter_0_avalon_slave_0_address -> arbiter_0:addr
	wire         mm_interconnect_0_arbiter_0_avalon_slave_0_read;                   // mm_interconnect_0:arbiter_0_avalon_slave_0_read -> arbiter_0:read
	wire         mm_interconnect_0_arbiter_0_avalon_slave_0_readdatavalid;          // arbiter_0:readack -> mm_interconnect_0:arbiter_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_arbiter_0_avalon_slave_0_write;                  // mm_interconnect_0:arbiter_0_avalon_slave_0_write -> arbiter_0:write
	wire   [7:0] mm_interconnect_0_arbiter_0_avalon_slave_0_writedata;              // mm_interconnect_0:arbiter_0_avalon_slave_0_writedata -> arbiter_0:din
	wire         mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_chipselect;  // mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_chipselect -> opencores_i2c:wb_cyc_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_readdata;    // opencores_i2c:wb_dat_o -> mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_readdata
	wire         mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_waitrequest; // opencores_i2c:wb_ack_o -> mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_waitrequest
	wire   [2:0] mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_address;     // mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_address -> opencores_i2c:wb_adr_i
	wire   [0:0] mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_byteenable;  // mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_byteenable -> opencores_i2c:wb_stb_i
	wire         mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_write;       // mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_write -> opencores_i2c:wb_we_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_writedata;   // mm_interconnect_0:opencores_i2c_bladerf_oc_i2c_master_writedata -> opencores_i2c:wb_dat_i
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                  // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;               // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;               // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                   // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                      // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                     // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                 // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_control_s1_chipselect;                           // mm_interconnect_0:control_s1_chipselect -> control:chipselect
	wire  [31:0] mm_interconnect_0_control_s1_readdata;                             // control:readdata -> mm_interconnect_0:control_s1_readdata
	wire   [2:0] mm_interconnect_0_control_s1_address;                              // mm_interconnect_0:control_s1_address -> control:address
	wire         mm_interconnect_0_control_s1_write;                                // mm_interconnect_0:control_s1_write -> control:write_n
	wire  [31:0] mm_interconnect_0_control_s1_writedata;                            // mm_interconnect_0:control_s1_writedata -> control:writedata
	wire         mm_interconnect_0_gpio_rffe_0_s1_chipselect;                       // mm_interconnect_0:gpio_rffe_0_s1_chipselect -> gpio_rffe_0:chipselect
	wire  [31:0] mm_interconnect_0_gpio_rffe_0_s1_readdata;                         // gpio_rffe_0:readdata -> mm_interconnect_0:gpio_rffe_0_s1_readdata
	wire   [2:0] mm_interconnect_0_gpio_rffe_0_s1_address;                          // mm_interconnect_0:gpio_rffe_0_s1_address -> gpio_rffe_0:address
	wire         mm_interconnect_0_gpio_rffe_0_s1_write;                            // mm_interconnect_0:gpio_rffe_0_s1_write -> gpio_rffe_0:write_n
	wire  [31:0] mm_interconnect_0_gpio_rffe_0_s1_writedata;                        // mm_interconnect_0:gpio_rffe_0_s1_writedata -> gpio_rffe_0:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                               // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                 // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [14:0] mm_interconnect_0_ram_s1_address;                                  // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                               // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                    // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                    // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_rx_trigger_ctl_s1_chipselect;                    // mm_interconnect_0:rx_trigger_ctl_s1_chipselect -> rx_trigger_ctl:chipselect
	wire  [31:0] mm_interconnect_0_rx_trigger_ctl_s1_readdata;                      // rx_trigger_ctl:readdata -> mm_interconnect_0:rx_trigger_ctl_s1_readdata
	wire   [2:0] mm_interconnect_0_rx_trigger_ctl_s1_address;                       // mm_interconnect_0:rx_trigger_ctl_s1_address -> rx_trigger_ctl:address
	wire         mm_interconnect_0_rx_trigger_ctl_s1_write;                         // mm_interconnect_0:rx_trigger_ctl_s1_write -> rx_trigger_ctl:write_n
	wire  [31:0] mm_interconnect_0_rx_trigger_ctl_s1_writedata;                     // mm_interconnect_0:rx_trigger_ctl_s1_writedata -> rx_trigger_ctl:writedata
	wire         mm_interconnect_0_tx_trigger_ctl_s1_chipselect;                    // mm_interconnect_0:tx_trigger_ctl_s1_chipselect -> tx_trigger_ctl:chipselect
	wire  [31:0] mm_interconnect_0_tx_trigger_ctl_s1_readdata;                      // tx_trigger_ctl:readdata -> mm_interconnect_0:tx_trigger_ctl_s1_readdata
	wire   [2:0] mm_interconnect_0_tx_trigger_ctl_s1_address;                       // mm_interconnect_0:tx_trigger_ctl_s1_address -> tx_trigger_ctl:address
	wire         mm_interconnect_0_tx_trigger_ctl_s1_write;                         // mm_interconnect_0:tx_trigger_ctl_s1_write -> tx_trigger_ctl:write_n
	wire  [31:0] mm_interconnect_0_tx_trigger_ctl_s1_writedata;                     // mm_interconnect_0:tx_trigger_ctl_s1_writedata -> tx_trigger_ctl:writedata
	wire         mm_interconnect_0_vctcxo_tamer_0_s1_chipselect;                    // mm_interconnect_0:vctcxo_tamer_0_s1_chipselect -> vctcxo_tamer_0:chipselect
	wire   [7:0] mm_interconnect_0_vctcxo_tamer_0_s1_readdata;                      // vctcxo_tamer_0:readdata -> mm_interconnect_0:vctcxo_tamer_0_s1_readdata
	wire   [7:0] mm_interconnect_0_vctcxo_tamer_0_s1_address;                       // mm_interconnect_0:vctcxo_tamer_0_s1_address -> vctcxo_tamer_0:address
	wire         mm_interconnect_0_vctcxo_tamer_0_s1_write;                         // mm_interconnect_0:vctcxo_tamer_0_s1_write -> vctcxo_tamer_0:write
	wire   [7:0] mm_interconnect_0_vctcxo_tamer_0_s1_writedata;                     // mm_interconnect_0:vctcxo_tamer_0_s1_writedata -> vctcxo_tamer_0:writedata
	wire         mm_interconnect_0_vctcxo_tamer_0_s1_clken;                         // mm_interconnect_0:vctcxo_tamer_0_s1_clken -> vctcxo_tamer_0:clken
	wire         mm_interconnect_0_xb_gpio_s1_chipselect;                           // mm_interconnect_0:xb_gpio_s1_chipselect -> xb_gpio:chipselect
	wire  [31:0] mm_interconnect_0_xb_gpio_s1_readdata;                             // xb_gpio:readdata -> mm_interconnect_0:xb_gpio_s1_readdata
	wire   [1:0] mm_interconnect_0_xb_gpio_s1_address;                              // mm_interconnect_0:xb_gpio_s1_address -> xb_gpio:address
	wire         mm_interconnect_0_xb_gpio_s1_write;                                // mm_interconnect_0:xb_gpio_s1_write -> xb_gpio:write_n
	wire  [31:0] mm_interconnect_0_xb_gpio_s1_writedata;                            // mm_interconnect_0:xb_gpio_s1_writedata -> xb_gpio:writedata
	wire         mm_interconnect_0_xb_gpio_dir_s1_chipselect;                       // mm_interconnect_0:xb_gpio_dir_s1_chipselect -> xb_gpio_dir:chipselect
	wire  [31:0] mm_interconnect_0_xb_gpio_dir_s1_readdata;                         // xb_gpio_dir:readdata -> mm_interconnect_0:xb_gpio_dir_s1_readdata
	wire   [1:0] mm_interconnect_0_xb_gpio_dir_s1_address;                          // mm_interconnect_0:xb_gpio_dir_s1_address -> xb_gpio_dir:address
	wire         mm_interconnect_0_xb_gpio_dir_s1_write;                            // mm_interconnect_0:xb_gpio_dir_s1_write -> xb_gpio_dir:write_n
	wire  [31:0] mm_interconnect_0_xb_gpio_dir_s1_writedata;                        // mm_interconnect_0:xb_gpio_dir_s1_writedata -> xb_gpio_dir:writedata
	wire  [15:0] mm_interconnect_0_axi_ad9361_0_s_axi_awaddr;                       // mm_interconnect_0:axi_ad9361_0_s_axi_awaddr -> axi_ad9361_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_ad9361_0_s_axi_bresp;                        // axi_ad9361_0:s_axi_bresp -> mm_interconnect_0:axi_ad9361_0_s_axi_bresp
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_arready;                      // axi_ad9361_0:s_axi_arready -> mm_interconnect_0:axi_ad9361_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_ad9361_0_s_axi_rdata;                        // axi_ad9361_0:s_axi_rdata -> mm_interconnect_0:axi_ad9361_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_ad9361_0_s_axi_wstrb;                        // mm_interconnect_0:axi_ad9361_0_s_axi_wstrb -> axi_ad9361_0:s_axi_wstrb
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_wready;                       // axi_ad9361_0:s_axi_wready -> mm_interconnect_0:axi_ad9361_0_s_axi_wready
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_awready;                      // axi_ad9361_0:s_axi_awready -> mm_interconnect_0:axi_ad9361_0_s_axi_awready
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_rready;                       // mm_interconnect_0:axi_ad9361_0_s_axi_rready -> axi_ad9361_0:s_axi_rready
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_bready;                       // mm_interconnect_0:axi_ad9361_0_s_axi_bready -> axi_ad9361_0:s_axi_bready
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_wvalid;                       // mm_interconnect_0:axi_ad9361_0_s_axi_wvalid -> axi_ad9361_0:s_axi_wvalid
	wire  [15:0] mm_interconnect_0_axi_ad9361_0_s_axi_araddr;                       // mm_interconnect_0:axi_ad9361_0_s_axi_araddr -> axi_ad9361_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_ad9361_0_s_axi_arprot;                       // mm_interconnect_0:axi_ad9361_0_s_axi_arprot -> axi_ad9361_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_ad9361_0_s_axi_rresp;                        // axi_ad9361_0:s_axi_rresp -> mm_interconnect_0:axi_ad9361_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_ad9361_0_s_axi_awprot;                       // mm_interconnect_0:axi_ad9361_0_s_axi_awprot -> axi_ad9361_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_ad9361_0_s_axi_wdata;                        // mm_interconnect_0:axi_ad9361_0_s_axi_wdata -> axi_ad9361_0:s_axi_wdata
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_arvalid;                      // mm_interconnect_0:axi_ad9361_0_s_axi_arvalid -> axi_ad9361_0:s_axi_arvalid
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_bvalid;                       // axi_ad9361_0:s_axi_bvalid -> mm_interconnect_0:axi_ad9361_0_s_axi_bvalid
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_awvalid;                      // mm_interconnect_0:axi_ad9361_0_s_axi_awvalid -> axi_ad9361_0:s_axi_awvalid
	wire         mm_interconnect_0_axi_ad9361_0_s_axi_rvalid;                       // axi_ad9361_0:s_axi_rvalid -> mm_interconnect_0:axi_ad9361_0_s_axi_rvalid
	wire         mm_interconnect_0_peripheral_spi_spi_control_port_chipselect;      // mm_interconnect_0:peripheral_spi_spi_control_port_chipselect -> peripheral_spi:spi_select
	wire  [15:0] mm_interconnect_0_peripheral_spi_spi_control_port_readdata;        // peripheral_spi:data_to_cpu -> mm_interconnect_0:peripheral_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_peripheral_spi_spi_control_port_address;         // mm_interconnect_0:peripheral_spi_spi_control_port_address -> peripheral_spi:mem_addr
	wire         mm_interconnect_0_peripheral_spi_spi_control_port_read;            // mm_interconnect_0:peripheral_spi_spi_control_port_read -> peripheral_spi:read_n
	wire         mm_interconnect_0_peripheral_spi_spi_control_port_write;           // mm_interconnect_0:peripheral_spi_spi_control_port_write -> peripheral_spi:write_n
	wire  [15:0] mm_interconnect_0_peripheral_spi_spi_control_port_writedata;       // mm_interconnect_0:peripheral_spi_spi_control_port_writedata -> peripheral_spi:data_from_cpu
	wire         mm_interconnect_0_rffe_spi_spi_control_port_chipselect;            // mm_interconnect_0:rffe_spi_spi_control_port_chipselect -> rffe_spi:spi_select
	wire  [15:0] mm_interconnect_0_rffe_spi_spi_control_port_readdata;              // rffe_spi:data_to_cpu -> mm_interconnect_0:rffe_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_rffe_spi_spi_control_port_address;               // mm_interconnect_0:rffe_spi_spi_control_port_address -> rffe_spi:mem_addr
	wire         mm_interconnect_0_rffe_spi_spi_control_port_read;                  // mm_interconnect_0:rffe_spi_spi_control_port_read -> rffe_spi:read_n
	wire         mm_interconnect_0_rffe_spi_spi_control_port_write;                 // mm_interconnect_0:rffe_spi_spi_control_port_write -> rffe_spi:write_n
	wire  [15:0] mm_interconnect_0_rffe_spi_spi_control_port_writedata;             // mm_interconnect_0:rffe_spi_spi_control_port_writedata -> rffe_spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                          // command_uart:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                          // arbiter_0:intr -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                          // opencores_i2c:wb_inta_o -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                          // rx_tamer:intr -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                          // wishbone_master_0:intr -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                          // tx_tamer:intr -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                          // gpio_rffe_0:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                          // peripheral_spi:irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                          // rffe_spi:irq -> irq_mapper:receiver9_irq
	wire  [31:0] nios2_irq_irq;                                                     // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [arbiter_0:reset, axi_ad9361_0:s_axi_aresetn, command_uart:reset, control:reset_n, gpio_rffe_0:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, opencores_i2c:wb_rst_i, peripheral_spi:reset_n, ram:reset, rffe_spi:reset_n, rst_translator:in_reset, rx_tamer:reset, rx_trigger_ctl:reset_n, tx_tamer:reset, tx_trigger_ctl:reset_n, vctcxo_tamer_0:reset, wishbone_master_0:reset, xb_gpio:reset_n, xb_gpio_dir:reset_n]
	wire         rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [nios2:reset_req, ram:reset_req, rst_translator:reset_req_in, vctcxo_tamer_0:reset_req]

	arbiter #(
		.N (2)
	) arbiter_0 (
		.addr    (mm_interconnect_0_arbiter_0_avalon_slave_0_address),       //   avalon_slave_0.address
		.din     (mm_interconnect_0_arbiter_0_avalon_slave_0_writedata),     //                 .writedata
		.dout    (mm_interconnect_0_arbiter_0_avalon_slave_0_readdata),      //                 .readdata
		.write   (mm_interconnect_0_arbiter_0_avalon_slave_0_write),         //                 .write
		.read    (mm_interconnect_0_arbiter_0_avalon_slave_0_read),          //                 .read
		.waitreq (mm_interconnect_0_arbiter_0_avalon_slave_0_waitrequest),   //                 .waitrequest
		.readack (mm_interconnect_0_arbiter_0_avalon_slave_0_readdatavalid), //                 .readdatavalid
		.reset   (rst_controller_reset_out_reset),                           //            reset.reset
		.request (arbiter_request),                                          //      conduit_end.request
		.granted (arbiter_granted),                                          //                 .granted
		.ack     (arbiter_ack),                                              //                 .ack
		.intr    (irq_mapper_receiver1_irq),                                 // interrupt_sender.irq
		.clock   (clk_clk)                                                   //       clock_sink.clk
	);

	axi_ad9361 #(
		.ID              (0),
		.DEVICE_TYPE     (0),
		.DAC_DDS_DISABLE (1)
	) axi_ad9361_0 (
		.s_axi_aclk     (clk_clk),                                      //     s_axi_clock.clk
		.s_axi_aresetn  (~rst_controller_reset_out_reset),              //     s_axi_reset.reset_n
		.s_axi_awvalid  (mm_interconnect_0_axi_ad9361_0_s_axi_awvalid), //           s_axi.awvalid
		.s_axi_awaddr   (mm_interconnect_0_axi_ad9361_0_s_axi_awaddr),  //                .awaddr
		.s_axi_awprot   (mm_interconnect_0_axi_ad9361_0_s_axi_awprot),  //                .awprot
		.s_axi_awready  (mm_interconnect_0_axi_ad9361_0_s_axi_awready), //                .awready
		.s_axi_wvalid   (mm_interconnect_0_axi_ad9361_0_s_axi_wvalid),  //                .wvalid
		.s_axi_wdata    (mm_interconnect_0_axi_ad9361_0_s_axi_wdata),   //                .wdata
		.s_axi_wstrb    (mm_interconnect_0_axi_ad9361_0_s_axi_wstrb),   //                .wstrb
		.s_axi_wready   (mm_interconnect_0_axi_ad9361_0_s_axi_wready),  //                .wready
		.s_axi_bvalid   (mm_interconnect_0_axi_ad9361_0_s_axi_bvalid),  //                .bvalid
		.s_axi_bresp    (mm_interconnect_0_axi_ad9361_0_s_axi_bresp),   //                .bresp
		.s_axi_bready   (mm_interconnect_0_axi_ad9361_0_s_axi_bready),  //                .bready
		.s_axi_arvalid  (mm_interconnect_0_axi_ad9361_0_s_axi_arvalid), //                .arvalid
		.s_axi_araddr   (mm_interconnect_0_axi_ad9361_0_s_axi_araddr),  //                .araddr
		.s_axi_arprot   (mm_interconnect_0_axi_ad9361_0_s_axi_arprot),  //                .arprot
		.s_axi_arready  (mm_interconnect_0_axi_ad9361_0_s_axi_arready), //                .arready
		.s_axi_rvalid   (mm_interconnect_0_axi_ad9361_0_s_axi_rvalid),  //                .rvalid
		.s_axi_rresp    (mm_interconnect_0_axi_ad9361_0_s_axi_rresp),   //                .rresp
		.s_axi_rdata    (mm_interconnect_0_axi_ad9361_0_s_axi_rdata),   //                .rdata
		.s_axi_rready   (mm_interconnect_0_axi_ad9361_0_s_axi_rready),  //                .rready
		.clk            (ad9361_data_clock_clk),                        //    device_clock.clk
		.rx_clk_in_p    (ad9361_device_if_rx_clk_in_p),                 //       device_if.rx_clk_in_p
		.rx_clk_in_n    (ad9361_device_if_rx_clk_in_n),                 //                .rx_clk_in_n
		.rx_frame_in_p  (ad9361_device_if_rx_frame_in_p),               //                .rx_frame_in_p
		.rx_frame_in_n  (ad9361_device_if_rx_frame_in_n),               //                .rx_frame_in_n
		.rx_data_in_p   (ad9361_device_if_rx_data_in_p),                //                .rx_data_in_p
		.rx_data_in_n   (ad9361_device_if_rx_data_in_n),                //                .rx_data_in_n
		.tx_clk_out_p   (ad9361_device_if_tx_clk_out_p),                //                .tx_clk_out_p
		.tx_clk_out_n   (ad9361_device_if_tx_clk_out_n),                //                .tx_clk_out_n
		.tx_frame_out_p (ad9361_device_if_tx_frame_out_p),              //                .tx_frame_out_p
		.tx_frame_out_n (ad9361_device_if_tx_frame_out_n),              //                .tx_frame_out_n
		.tx_data_out_p  (ad9361_device_if_tx_data_out_p),               //                .tx_data_out_p
		.tx_data_out_n  (ad9361_device_if_tx_data_out_n),               //                .tx_data_out_n
		.dac_sync_in    (ad9361_dac_sync_in_sync),                      //  if_dac_sync_in.sync
		.dac_sync_out   (ad9361_dac_sync_out_sync),                     // if_dac_sync_out.sync
		.l_clk          (ad9361_data_clock_clk),                        //        if_l_clk.clk
		.rst            (ad9361_data_reset_reset),                      //          if_rst.reset
		.adc_enable_i0  (ad9361_adc_i0_enable),                         //    fifo_ch_0_in.enable
		.adc_valid_i0   (ad9361_adc_i0_valid),                          //                .valid
		.adc_data_i0    (ad9361_adc_i0_data),                           //                .data
		.adc_enable_q0  (ad9361_adc_q0_enable),                         //    fifo_ch_1_in.enable
		.adc_valid_q0   (ad9361_adc_q0_valid),                          //                .valid
		.adc_data_q0    (ad9361_adc_q0_data),                           //                .data
		.adc_enable_i1  (ad9361_adc_i1_enable),                         //    fifo_ch_2_in.enable
		.adc_valid_i1   (ad9361_adc_i1_valid),                          //                .valid
		.adc_data_i1    (ad9361_adc_i1_data),                           //                .data
		.adc_enable_q1  (ad9361_adc_q1_enable),                         //    fifo_ch_3_in.enable
		.adc_valid_q1   (ad9361_adc_q1_valid),                          //                .valid
		.adc_data_q1    (ad9361_adc_q1_data),                           //                .data
		.adc_dovf       (ad9361_adc_overflow_ovf),                      //     if_adc_dovf.ovf
		.adc_dunf       (ad9361_adc_underflow_unf),                     //     if_adc_dunf.unf
		.dac_enable_i0  (ad9361_dac_i0_enable),                         //   fifo_ch_0_out.enable
		.dac_valid_i0   (ad9361_dac_i0_valid),                          //                .valid
		.dac_data_i0    (ad9361_dac_i0_data),                           //                .data
		.dac_enable_q0  (ad9361_dac_q0_enable),                         //   fifo_ch_1_out.enable
		.dac_valid_q0   (ad9361_dac_q0_valid),                          //                .valid
		.dac_data_q0    (ad9361_dac_q0_data),                           //                .data
		.dac_enable_i1  (ad9361_dac_i1_enable),                         //   fifo_ch_2_out.enable
		.dac_valid_i1   (ad9361_dac_i1_valid),                          //                .valid
		.dac_data_i1    (ad9361_dac_i1_data),                           //                .data
		.dac_enable_q1  (ad9361_dac_q1_enable),                         //   fifo_ch_3_out.enable
		.dac_valid_q1   (ad9361_dac_q1_valid),                          //                .valid
		.dac_data_q1    (ad9361_dac_q1_data),                           //                .data
		.dac_dovf       (ad9361_dac_overflow_ovf),                      //     if_dac_dovf.ovf
		.dac_dunf       (ad9361_dac_underflow_unf),                     //     if_dac_dunf.unf
		.delay_clk      (clk_clk)                                       //     delay_clock.clk
	);

	command_uart command_uart (
		.reset      (rst_controller_reset_out_reset),                            //        reset.reset
		.rs232_sin  (command_serial_in),                                         //        rs232.serial_in
		.rs232_sout (command_serial_out),                                        //             .serial_out
		.irq        (irq_mapper_receiver0_irq),                                  //    interrupt.irq
		.clock      (clk_clk),                                                   //        clock.clk
		.addr       (mm_interconnect_0_command_uart_avalon_slave_address),       // avalon_slave.address
		.dout       (mm_interconnect_0_command_uart_avalon_slave_readdata),      //             .readdata
		.din        (mm_interconnect_0_command_uart_avalon_slave_writedata),     //             .writedata
		.read       (mm_interconnect_0_command_uart_avalon_slave_read),          //             .read
		.write      (mm_interconnect_0_command_uart_avalon_slave_write),         //             .write
		.readack    (mm_interconnect_0_command_uart_avalon_slave_readdatavalid), //             .readdatavalid
		.waitreq    (mm_interconnect_0_command_uart_avalon_slave_waitrequest)    //             .waitrequest
	);

	nios_system_control control (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_control_s1_readdata),   //                    .readdata
		.in_port    (gpio_in_port),                            // external_connection.export
		.out_port   (gpio_out_port)                            //                    .export
	);

	nios_system_gpio_rffe_0 gpio_rffe_0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_gpio_rffe_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_rffe_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_rffe_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_rffe_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_rffe_0_s1_readdata),   //                    .readdata
		.in_port    (gpio_rffe_0_in_port),                         // external_connection.export
		.out_port   (gpio_rffe_0_out_port),                        //                    .export
		.irq        (irq_mapper_receiver6_irq)                     //                 irq.irq
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver7_irq)                                   //               irq.irq
	);

	nios_system_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	i2c_master_top #(
		.ARST_LVL (1)
	) opencores_i2c (
		.wb_clk_i     (clk_clk),                                                           //            clock_sink.clk
		.wb_rst_i     (rst_controller_reset_out_reset),                                    //            reset_sink.reset
		.scl_pad_o    (oc_i2c_scl_pad_o),                                                  //           conduit_end.scl_pad_o
		.scl_padoen_o (oc_i2c_scl_padoen_o),                                               //                      .scl_padoen_o
		.sda_pad_i    (oc_i2c_sda_pad_i),                                                  //                      .sda_pad_i
		.sda_pad_o    (oc_i2c_sda_pad_o),                                                  //                      .sda_pad_o
		.sda_padoen_o (oc_i2c_sda_padoen_o),                                               //                      .sda_padoen_o
		.arst_i       (oc_i2c_arst_i),                                                     //                      .arst_i
		.scl_pad_i    (oc_i2c_scl_pad_i),                                                  //                      .scl_pad_i
		.wb_inta_o    (irq_mapper_receiver2_irq),                                          //      interrupt_sender.irq
		.wb_dat_i     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_writedata),   // bladerf_oc_i2c_master.writedata
		.wb_dat_o     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_readdata),    //                      .readdata
		.wb_we_i      (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_write),       //                      .write
		.wb_stb_i     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_byteenable),  //                      .byteenable
		.wb_cyc_i     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_chipselect),  //                      .chipselect
		.wb_ack_o     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_waitrequest), //                      .waitrequest_n
		.wb_adr_i     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_address)      //                      .address
	);

	nios_system_peripheral_spi peripheral_spi (
		.clk           (clk_clk),                                                      //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                              //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_peripheral_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_peripheral_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_peripheral_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_peripheral_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_peripheral_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_peripheral_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver8_irq),                                     //              irq.irq
		.MISO          (dac_MISO),                                                     //         external.export
		.MOSI          (dac_MOSI),                                                     //                 .export
		.SCLK          (dac_SCLK),                                                     //                 .export
		.SS_n          (dac_SS_n)                                                      //                 .export
	);

	nios_system_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	nios_system_rffe_spi rffe_spi (
		.clk           (clk_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_rffe_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_rffe_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_rffe_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_rffe_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_rffe_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_rffe_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver9_irq),                               //              irq.irq
		.MISO          (spi_MISO),                                               //         external.export
		.MOSI          (spi_MOSI),                                               //                 .export
		.SCLK          (spi_SCLK),                                               //                 .export
		.SS_n          (spi_SS_n)                                                //                 .export
	);

	time_tamer rx_tamer (
		.reset       (rst_controller_reset_out_reset),                          //            reset.reset
		.din         (mm_interconnect_0_rx_tamer_avalon_slave_0_writedata),     //   avalon_slave_0.writedata
		.dout        (mm_interconnect_0_rx_tamer_avalon_slave_0_readdata),      //                 .readdata
		.write       (mm_interconnect_0_rx_tamer_avalon_slave_0_write),         //                 .write
		.read        (mm_interconnect_0_rx_tamer_avalon_slave_0_read),          //                 .read
		.waitreq     (mm_interconnect_0_rx_tamer_avalon_slave_0_waitrequest),   //                 .waitrequest
		.readack     (mm_interconnect_0_rx_tamer_avalon_slave_0_readdatavalid), //                 .readdatavalid
		.addr        (mm_interconnect_0_rx_tamer_avalon_slave_0_address),       //                 .address
		.clock       (clk_clk),                                                 //       clock_sink.clk
		.intr        (irq_mapper_receiver3_irq),                                // interrupt_sender.irq
		.ts_sync_in  (rx_tamer_ts_sync_in),                                     //      conduit_end.ts_sync_in
		.ts_sync_out (rx_tamer_ts_sync_out),                                    //                 .ts_sync_out
		.ts_pps      (rx_tamer_ts_pps),                                         //                 .ts_pps
		.ts_clock    (rx_tamer_ts_clock),                                       //                 .ts_clock
		.ts_reset    (rx_tamer_ts_reset),                                       //                 .ts_reset
		.ts_time     (rx_tamer_ts_time)                                         //                 .ts_time
	);

	nios_system_rx_trigger_ctl rx_trigger_ctl (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_rx_trigger_ctl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rx_trigger_ctl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rx_trigger_ctl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rx_trigger_ctl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rx_trigger_ctl_s1_readdata),   //                    .readdata
		.in_port    (rx_trigger_ctl_in_port),                         // external_connection.export
		.out_port   (rx_trigger_ctl_out_port)                         //                    .export
	);

	time_tamer tx_tamer (
		.reset       (rst_controller_reset_out_reset),                          //            reset.reset
		.din         (mm_interconnect_0_tx_tamer_avalon_slave_0_writedata),     //   avalon_slave_0.writedata
		.dout        (mm_interconnect_0_tx_tamer_avalon_slave_0_readdata),      //                 .readdata
		.write       (mm_interconnect_0_tx_tamer_avalon_slave_0_write),         //                 .write
		.read        (mm_interconnect_0_tx_tamer_avalon_slave_0_read),          //                 .read
		.waitreq     (mm_interconnect_0_tx_tamer_avalon_slave_0_waitrequest),   //                 .waitrequest
		.readack     (mm_interconnect_0_tx_tamer_avalon_slave_0_readdatavalid), //                 .readdatavalid
		.addr        (mm_interconnect_0_tx_tamer_avalon_slave_0_address),       //                 .address
		.clock       (clk_clk),                                                 //       clock_sink.clk
		.intr        (irq_mapper_receiver5_irq),                                // interrupt_sender.irq
		.ts_sync_in  (tx_tamer_ts_sync_in),                                     //      conduit_end.ts_sync_in
		.ts_sync_out (tx_tamer_ts_sync_out),                                    //                 .ts_sync_out
		.ts_pps      (tx_tamer_ts_pps),                                         //                 .ts_pps
		.ts_clock    (tx_tamer_ts_clock),                                       //                 .ts_clock
		.ts_reset    (tx_tamer_ts_reset),                                       //                 .ts_reset
		.ts_time     (tx_tamer_ts_time)                                         //                 .ts_time
	);

	nios_system_rx_trigger_ctl tx_trigger_ctl (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_tx_trigger_ctl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tx_trigger_ctl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tx_trigger_ctl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tx_trigger_ctl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tx_trigger_ctl_s1_readdata),   //                    .readdata
		.in_port    (tx_trigger_ctl_in_port),                         // external_connection.export
		.out_port   (tx_trigger_ctl_out_port)                         //                    .export
	);

	nios_system_vctcxo_tamer_0 vctcxo_tamer_0 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_vctcxo_tamer_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_vctcxo_tamer_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_vctcxo_tamer_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_vctcxo_tamer_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_vctcxo_tamer_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_vctcxo_tamer_0_s1_writedata),  //       .writedata
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	wishbone_master #(
		.ADDR_BITS (32),
		.DATA_BITS (32)
	) wishbone_master_0 (
		.addr     (mm_interconnect_0_wishbone_master_0_avalon_slave_0_address),       //   avalon_slave_0.address
		.din      (mm_interconnect_0_wishbone_master_0_avalon_slave_0_writedata),     //                 .writedata
		.dout     (mm_interconnect_0_wishbone_master_0_avalon_slave_0_readdata),      //                 .readdata
		.write    (mm_interconnect_0_wishbone_master_0_avalon_slave_0_write),         //                 .write
		.read     (mm_interconnect_0_wishbone_master_0_avalon_slave_0_read),          //                 .read
		.waitreq  (mm_interconnect_0_wishbone_master_0_avalon_slave_0_waitrequest),   //                 .waitrequest
		.readack  (mm_interconnect_0_wishbone_master_0_avalon_slave_0_readdatavalid), //                 .readdatavalid
		.reset    (rst_controller_reset_out_reset),                                   //            reset.reset
		.wb_clk_i (wbm_wb_clk_i),                                                     //      conduit_end.wb_clk_i
		.wb_rst_i (wbm_wb_rst_i),                                                     //                 .wb_rst_i
		.wb_adr_o (wbm_wb_adr_o),                                                     //                 .wb_adr_o
		.wb_dat_o (wbm_wb_dat_o),                                                     //                 .wb_dat_o
		.wb_dat_i (wbm_wb_dat_i),                                                     //                 .wb_dat_i
		.wb_we_o  (wbm_wb_we_o),                                                      //                 .wb_we_o
		.wb_sel_o (wbm_wb_sel_o),                                                     //                 .wb_sel_o
		.wb_stb_o (wbm_wb_stb_o),                                                     //                 .wb_stb_o
		.wb_ack_i (wbm_wb_ack_i),                                                     //                 .wb_ack_i
		.wb_cyc_o (wbm_wb_cyc_o),                                                     //                 .wb_cyc_o
		.intr     (irq_mapper_receiver4_irq),                                         // interrupt_sender.irq
		.clock    (clk_clk)                                                           //       clock_sink.clk
	);

	nios_system_xb_gpio xb_gpio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_xb_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_xb_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_xb_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_xb_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_xb_gpio_s1_readdata),   //                    .readdata
		.in_port    (xb_gpio_in_port),                         // external_connection.export
		.out_port   (xb_gpio_out_port)                         //                    .export
	);

	nios_system_xb_gpio_dir xb_gpio_dir (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_xb_gpio_dir_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_xb_gpio_dir_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_xb_gpio_dir_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_xb_gpio_dir_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_xb_gpio_dir_s1_readdata),   //                    .readdata
		.out_port   (xb_gpio_dir_export)                           // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.axi_ad9361_0_s_axi_awaddr                       (mm_interconnect_0_axi_ad9361_0_s_axi_awaddr),                        //                  axi_ad9361_0_s_axi.awaddr
		.axi_ad9361_0_s_axi_awprot                       (mm_interconnect_0_axi_ad9361_0_s_axi_awprot),                        //                                    .awprot
		.axi_ad9361_0_s_axi_awvalid                      (mm_interconnect_0_axi_ad9361_0_s_axi_awvalid),                       //                                    .awvalid
		.axi_ad9361_0_s_axi_awready                      (mm_interconnect_0_axi_ad9361_0_s_axi_awready),                       //                                    .awready
		.axi_ad9361_0_s_axi_wdata                        (mm_interconnect_0_axi_ad9361_0_s_axi_wdata),                         //                                    .wdata
		.axi_ad9361_0_s_axi_wstrb                        (mm_interconnect_0_axi_ad9361_0_s_axi_wstrb),                         //                                    .wstrb
		.axi_ad9361_0_s_axi_wvalid                       (mm_interconnect_0_axi_ad9361_0_s_axi_wvalid),                        //                                    .wvalid
		.axi_ad9361_0_s_axi_wready                       (mm_interconnect_0_axi_ad9361_0_s_axi_wready),                        //                                    .wready
		.axi_ad9361_0_s_axi_bresp                        (mm_interconnect_0_axi_ad9361_0_s_axi_bresp),                         //                                    .bresp
		.axi_ad9361_0_s_axi_bvalid                       (mm_interconnect_0_axi_ad9361_0_s_axi_bvalid),                        //                                    .bvalid
		.axi_ad9361_0_s_axi_bready                       (mm_interconnect_0_axi_ad9361_0_s_axi_bready),                        //                                    .bready
		.axi_ad9361_0_s_axi_araddr                       (mm_interconnect_0_axi_ad9361_0_s_axi_araddr),                        //                                    .araddr
		.axi_ad9361_0_s_axi_arprot                       (mm_interconnect_0_axi_ad9361_0_s_axi_arprot),                        //                                    .arprot
		.axi_ad9361_0_s_axi_arvalid                      (mm_interconnect_0_axi_ad9361_0_s_axi_arvalid),                       //                                    .arvalid
		.axi_ad9361_0_s_axi_arready                      (mm_interconnect_0_axi_ad9361_0_s_axi_arready),                       //                                    .arready
		.axi_ad9361_0_s_axi_rdata                        (mm_interconnect_0_axi_ad9361_0_s_axi_rdata),                         //                                    .rdata
		.axi_ad9361_0_s_axi_rresp                        (mm_interconnect_0_axi_ad9361_0_s_axi_rresp),                         //                                    .rresp
		.axi_ad9361_0_s_axi_rvalid                       (mm_interconnect_0_axi_ad9361_0_s_axi_rvalid),                        //                                    .rvalid
		.axi_ad9361_0_s_axi_rready                       (mm_interconnect_0_axi_ad9361_0_s_axi_rready),                        //                                    .rready
		.system_clock_clk_clk                            (clk_clk),                                                            //                    system_clock_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                     //   nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                       (nios2_data_master_address),                                          //                   nios2_data_master.address
		.nios2_data_master_waitrequest                   (nios2_data_master_waitrequest),                                      //                                    .waitrequest
		.nios2_data_master_byteenable                    (nios2_data_master_byteenable),                                       //                                    .byteenable
		.nios2_data_master_read                          (nios2_data_master_read),                                             //                                    .read
		.nios2_data_master_readdata                      (nios2_data_master_readdata),                                         //                                    .readdata
		.nios2_data_master_write                         (nios2_data_master_write),                                            //                                    .write
		.nios2_data_master_writedata                     (nios2_data_master_writedata),                                        //                                    .writedata
		.nios2_data_master_debugaccess                   (nios2_data_master_debugaccess),                                      //                                    .debugaccess
		.nios2_instruction_master_address                (nios2_instruction_master_address),                                   //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest            (nios2_instruction_master_waitrequest),                               //                                    .waitrequest
		.nios2_instruction_master_read                   (nios2_instruction_master_read),                                      //                                    .read
		.nios2_instruction_master_readdata               (nios2_instruction_master_readdata),                                  //                                    .readdata
		.arbiter_0_avalon_slave_0_address                (mm_interconnect_0_arbiter_0_avalon_slave_0_address),                 //            arbiter_0_avalon_slave_0.address
		.arbiter_0_avalon_slave_0_write                  (mm_interconnect_0_arbiter_0_avalon_slave_0_write),                   //                                    .write
		.arbiter_0_avalon_slave_0_read                   (mm_interconnect_0_arbiter_0_avalon_slave_0_read),                    //                                    .read
		.arbiter_0_avalon_slave_0_readdata               (mm_interconnect_0_arbiter_0_avalon_slave_0_readdata),                //                                    .readdata
		.arbiter_0_avalon_slave_0_writedata              (mm_interconnect_0_arbiter_0_avalon_slave_0_writedata),               //                                    .writedata
		.arbiter_0_avalon_slave_0_readdatavalid          (mm_interconnect_0_arbiter_0_avalon_slave_0_readdatavalid),           //                                    .readdatavalid
		.arbiter_0_avalon_slave_0_waitrequest            (mm_interconnect_0_arbiter_0_avalon_slave_0_waitrequest),             //                                    .waitrequest
		.command_uart_avalon_slave_address               (mm_interconnect_0_command_uart_avalon_slave_address),                //           command_uart_avalon_slave.address
		.command_uart_avalon_slave_write                 (mm_interconnect_0_command_uart_avalon_slave_write),                  //                                    .write
		.command_uart_avalon_slave_read                  (mm_interconnect_0_command_uart_avalon_slave_read),                   //                                    .read
		.command_uart_avalon_slave_readdata              (mm_interconnect_0_command_uart_avalon_slave_readdata),               //                                    .readdata
		.command_uart_avalon_slave_writedata             (mm_interconnect_0_command_uart_avalon_slave_writedata),              //                                    .writedata
		.command_uart_avalon_slave_readdatavalid         (mm_interconnect_0_command_uart_avalon_slave_readdatavalid),          //                                    .readdatavalid
		.command_uart_avalon_slave_waitrequest           (mm_interconnect_0_command_uart_avalon_slave_waitrequest),            //                                    .waitrequest
		.control_s1_address                              (mm_interconnect_0_control_s1_address),                               //                          control_s1.address
		.control_s1_write                                (mm_interconnect_0_control_s1_write),                                 //                                    .write
		.control_s1_readdata                             (mm_interconnect_0_control_s1_readdata),                              //                                    .readdata
		.control_s1_writedata                            (mm_interconnect_0_control_s1_writedata),                             //                                    .writedata
		.control_s1_chipselect                           (mm_interconnect_0_control_s1_chipselect),                            //                                    .chipselect
		.gpio_rffe_0_s1_address                          (mm_interconnect_0_gpio_rffe_0_s1_address),                           //                      gpio_rffe_0_s1.address
		.gpio_rffe_0_s1_write                            (mm_interconnect_0_gpio_rffe_0_s1_write),                             //                                    .write
		.gpio_rffe_0_s1_readdata                         (mm_interconnect_0_gpio_rffe_0_s1_readdata),                          //                                    .readdata
		.gpio_rffe_0_s1_writedata                        (mm_interconnect_0_gpio_rffe_0_s1_writedata),                         //                                    .writedata
		.gpio_rffe_0_s1_chipselect                       (mm_interconnect_0_gpio_rffe_0_s1_chipselect),                        //                                    .chipselect
		.jtag_uart_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                    .write
		.jtag_uart_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                    .chipselect
		.nios2_debug_mem_slave_address                   (mm_interconnect_0_nios2_debug_mem_slave_address),                    //               nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                     (mm_interconnect_0_nios2_debug_mem_slave_write),                      //                                    .write
		.nios2_debug_mem_slave_read                      (mm_interconnect_0_nios2_debug_mem_slave_read),                       //                                    .read
		.nios2_debug_mem_slave_readdata                  (mm_interconnect_0_nios2_debug_mem_slave_readdata),                   //                                    .readdata
		.nios2_debug_mem_slave_writedata                 (mm_interconnect_0_nios2_debug_mem_slave_writedata),                  //                                    .writedata
		.nios2_debug_mem_slave_byteenable                (mm_interconnect_0_nios2_debug_mem_slave_byteenable),                 //                                    .byteenable
		.nios2_debug_mem_slave_waitrequest               (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),                //                                    .waitrequest
		.nios2_debug_mem_slave_debugaccess               (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),                //                                    .debugaccess
		.opencores_i2c_bladerf_oc_i2c_master_address     (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_address),      // opencores_i2c_bladerf_oc_i2c_master.address
		.opencores_i2c_bladerf_oc_i2c_master_write       (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_write),        //                                    .write
		.opencores_i2c_bladerf_oc_i2c_master_readdata    (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_readdata),     //                                    .readdata
		.opencores_i2c_bladerf_oc_i2c_master_writedata   (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_writedata),    //                                    .writedata
		.opencores_i2c_bladerf_oc_i2c_master_byteenable  (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_byteenable),   //                                    .byteenable
		.opencores_i2c_bladerf_oc_i2c_master_waitrequest (~mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_waitrequest), //                                    .waitrequest
		.opencores_i2c_bladerf_oc_i2c_master_chipselect  (mm_interconnect_0_opencores_i2c_bladerf_oc_i2c_master_chipselect),   //                                    .chipselect
		.peripheral_spi_spi_control_port_address         (mm_interconnect_0_peripheral_spi_spi_control_port_address),          //     peripheral_spi_spi_control_port.address
		.peripheral_spi_spi_control_port_write           (mm_interconnect_0_peripheral_spi_spi_control_port_write),            //                                    .write
		.peripheral_spi_spi_control_port_read            (mm_interconnect_0_peripheral_spi_spi_control_port_read),             //                                    .read
		.peripheral_spi_spi_control_port_readdata        (mm_interconnect_0_peripheral_spi_spi_control_port_readdata),         //                                    .readdata
		.peripheral_spi_spi_control_port_writedata       (mm_interconnect_0_peripheral_spi_spi_control_port_writedata),        //                                    .writedata
		.peripheral_spi_spi_control_port_chipselect      (mm_interconnect_0_peripheral_spi_spi_control_port_chipselect),       //                                    .chipselect
		.ram_s1_address                                  (mm_interconnect_0_ram_s1_address),                                   //                              ram_s1.address
		.ram_s1_write                                    (mm_interconnect_0_ram_s1_write),                                     //                                    .write
		.ram_s1_readdata                                 (mm_interconnect_0_ram_s1_readdata),                                  //                                    .readdata
		.ram_s1_writedata                                (mm_interconnect_0_ram_s1_writedata),                                 //                                    .writedata
		.ram_s1_byteenable                               (mm_interconnect_0_ram_s1_byteenable),                                //                                    .byteenable
		.ram_s1_chipselect                               (mm_interconnect_0_ram_s1_chipselect),                                //                                    .chipselect
		.ram_s1_clken                                    (mm_interconnect_0_ram_s1_clken),                                     //                                    .clken
		.rffe_spi_spi_control_port_address               (mm_interconnect_0_rffe_spi_spi_control_port_address),                //           rffe_spi_spi_control_port.address
		.rffe_spi_spi_control_port_write                 (mm_interconnect_0_rffe_spi_spi_control_port_write),                  //                                    .write
		.rffe_spi_spi_control_port_read                  (mm_interconnect_0_rffe_spi_spi_control_port_read),                   //                                    .read
		.rffe_spi_spi_control_port_readdata              (mm_interconnect_0_rffe_spi_spi_control_port_readdata),               //                                    .readdata
		.rffe_spi_spi_control_port_writedata             (mm_interconnect_0_rffe_spi_spi_control_port_writedata),              //                                    .writedata
		.rffe_spi_spi_control_port_chipselect            (mm_interconnect_0_rffe_spi_spi_control_port_chipselect),             //                                    .chipselect
		.rx_tamer_avalon_slave_0_address                 (mm_interconnect_0_rx_tamer_avalon_slave_0_address),                  //             rx_tamer_avalon_slave_0.address
		.rx_tamer_avalon_slave_0_write                   (mm_interconnect_0_rx_tamer_avalon_slave_0_write),                    //                                    .write
		.rx_tamer_avalon_slave_0_read                    (mm_interconnect_0_rx_tamer_avalon_slave_0_read),                     //                                    .read
		.rx_tamer_avalon_slave_0_readdata                (mm_interconnect_0_rx_tamer_avalon_slave_0_readdata),                 //                                    .readdata
		.rx_tamer_avalon_slave_0_writedata               (mm_interconnect_0_rx_tamer_avalon_slave_0_writedata),                //                                    .writedata
		.rx_tamer_avalon_slave_0_readdatavalid           (mm_interconnect_0_rx_tamer_avalon_slave_0_readdatavalid),            //                                    .readdatavalid
		.rx_tamer_avalon_slave_0_waitrequest             (mm_interconnect_0_rx_tamer_avalon_slave_0_waitrequest),              //                                    .waitrequest
		.rx_trigger_ctl_s1_address                       (mm_interconnect_0_rx_trigger_ctl_s1_address),                        //                   rx_trigger_ctl_s1.address
		.rx_trigger_ctl_s1_write                         (mm_interconnect_0_rx_trigger_ctl_s1_write),                          //                                    .write
		.rx_trigger_ctl_s1_readdata                      (mm_interconnect_0_rx_trigger_ctl_s1_readdata),                       //                                    .readdata
		.rx_trigger_ctl_s1_writedata                     (mm_interconnect_0_rx_trigger_ctl_s1_writedata),                      //                                    .writedata
		.rx_trigger_ctl_s1_chipselect                    (mm_interconnect_0_rx_trigger_ctl_s1_chipselect),                     //                                    .chipselect
		.tx_tamer_avalon_slave_0_address                 (mm_interconnect_0_tx_tamer_avalon_slave_0_address),                  //             tx_tamer_avalon_slave_0.address
		.tx_tamer_avalon_slave_0_write                   (mm_interconnect_0_tx_tamer_avalon_slave_0_write),                    //                                    .write
		.tx_tamer_avalon_slave_0_read                    (mm_interconnect_0_tx_tamer_avalon_slave_0_read),                     //                                    .read
		.tx_tamer_avalon_slave_0_readdata                (mm_interconnect_0_tx_tamer_avalon_slave_0_readdata),                 //                                    .readdata
		.tx_tamer_avalon_slave_0_writedata               (mm_interconnect_0_tx_tamer_avalon_slave_0_writedata),                //                                    .writedata
		.tx_tamer_avalon_slave_0_readdatavalid           (mm_interconnect_0_tx_tamer_avalon_slave_0_readdatavalid),            //                                    .readdatavalid
		.tx_tamer_avalon_slave_0_waitrequest             (mm_interconnect_0_tx_tamer_avalon_slave_0_waitrequest),              //                                    .waitrequest
		.tx_trigger_ctl_s1_address                       (mm_interconnect_0_tx_trigger_ctl_s1_address),                        //                   tx_trigger_ctl_s1.address
		.tx_trigger_ctl_s1_write                         (mm_interconnect_0_tx_trigger_ctl_s1_write),                          //                                    .write
		.tx_trigger_ctl_s1_readdata                      (mm_interconnect_0_tx_trigger_ctl_s1_readdata),                       //                                    .readdata
		.tx_trigger_ctl_s1_writedata                     (mm_interconnect_0_tx_trigger_ctl_s1_writedata),                      //                                    .writedata
		.tx_trigger_ctl_s1_chipselect                    (mm_interconnect_0_tx_trigger_ctl_s1_chipselect),                     //                                    .chipselect
		.vctcxo_tamer_0_s1_address                       (mm_interconnect_0_vctcxo_tamer_0_s1_address),                        //                   vctcxo_tamer_0_s1.address
		.vctcxo_tamer_0_s1_write                         (mm_interconnect_0_vctcxo_tamer_0_s1_write),                          //                                    .write
		.vctcxo_tamer_0_s1_readdata                      (mm_interconnect_0_vctcxo_tamer_0_s1_readdata),                       //                                    .readdata
		.vctcxo_tamer_0_s1_writedata                     (mm_interconnect_0_vctcxo_tamer_0_s1_writedata),                      //                                    .writedata
		.vctcxo_tamer_0_s1_chipselect                    (mm_interconnect_0_vctcxo_tamer_0_s1_chipselect),                     //                                    .chipselect
		.vctcxo_tamer_0_s1_clken                         (mm_interconnect_0_vctcxo_tamer_0_s1_clken),                          //                                    .clken
		.wishbone_master_0_avalon_slave_0_address        (mm_interconnect_0_wishbone_master_0_avalon_slave_0_address),         //    wishbone_master_0_avalon_slave_0.address
		.wishbone_master_0_avalon_slave_0_write          (mm_interconnect_0_wishbone_master_0_avalon_slave_0_write),           //                                    .write
		.wishbone_master_0_avalon_slave_0_read           (mm_interconnect_0_wishbone_master_0_avalon_slave_0_read),            //                                    .read
		.wishbone_master_0_avalon_slave_0_readdata       (mm_interconnect_0_wishbone_master_0_avalon_slave_0_readdata),        //                                    .readdata
		.wishbone_master_0_avalon_slave_0_writedata      (mm_interconnect_0_wishbone_master_0_avalon_slave_0_writedata),       //                                    .writedata
		.wishbone_master_0_avalon_slave_0_readdatavalid  (mm_interconnect_0_wishbone_master_0_avalon_slave_0_readdatavalid),   //                                    .readdatavalid
		.wishbone_master_0_avalon_slave_0_waitrequest    (mm_interconnect_0_wishbone_master_0_avalon_slave_0_waitrequest),     //                                    .waitrequest
		.xb_gpio_s1_address                              (mm_interconnect_0_xb_gpio_s1_address),                               //                          xb_gpio_s1.address
		.xb_gpio_s1_write                                (mm_interconnect_0_xb_gpio_s1_write),                                 //                                    .write
		.xb_gpio_s1_readdata                             (mm_interconnect_0_xb_gpio_s1_readdata),                              //                                    .readdata
		.xb_gpio_s1_writedata                            (mm_interconnect_0_xb_gpio_s1_writedata),                             //                                    .writedata
		.xb_gpio_s1_chipselect                           (mm_interconnect_0_xb_gpio_s1_chipselect),                            //                                    .chipselect
		.xb_gpio_dir_s1_address                          (mm_interconnect_0_xb_gpio_dir_s1_address),                           //                      xb_gpio_dir_s1.address
		.xb_gpio_dir_s1_write                            (mm_interconnect_0_xb_gpio_dir_s1_write),                             //                                    .write
		.xb_gpio_dir_s1_readdata                         (mm_interconnect_0_xb_gpio_dir_s1_readdata),                          //                                    .readdata
		.xb_gpio_dir_s1_writedata                        (mm_interconnect_0_xb_gpio_dir_s1_writedata),                         //                                    .writedata
		.xb_gpio_dir_s1_chipselect                       (mm_interconnect_0_xb_gpio_dir_s1_chipselect)                         //                                    .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq),       // receiver9.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
