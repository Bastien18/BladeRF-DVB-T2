��/  �-�߰B�P��ي�m���+8�KS�����B������+�rz���C�
c�_����b-�����<�k
�9:K��J�g��$�u�m��	����l�i��,��F�.��[6�ө��_X��w��Mi���]�R��K��f�[c�Se�}{r`����C������U@G[l�Gݹ��W{���ȑ�����	e����Б�䷒5k,���*�'oP�'Fz�q�3�z���XۉERl�"�t�Eޠ��f+�yD�]�X0/���7��l��'��YŌ�=��1���^�9|�r�w�8�#gXN	��@����A�,��A�𞪐j�`XؾG8�S�F�䏬����tZ1I��Z�㓬�c�y}j� ��c~��K��k�\����n�-��[� ���4�"��B�=~����D��-�R���^Ƣ$����Y++�WL2t4?��>��=����,��.��Tt/]x���!;�\��[�x�e\6��،����ج8:۲ߊ�*.ѷ�E��\:Ϸ���1�x*�e�}��0�0��a�5L<���ݮ
r���\.q�6�����Ӝ������9����+�HEh�aE��l�O��:Xұ�U6n�Df ��y�J��� �ij�\�ΧU�א�)+)磳vzV��	�&�Lď�$�n�9@�:t:���O)g,K�[u��yΟ���0�A�&^������
D{�	򜴉�@� I#��e�� ���p3&@��o����]�D�	�(]���%���z�Q��=R���?�y��'��Kdܵ%Ԅ��_@�"zT�>܃n�~��Q�9{��$y�:{��b�؏��`�$�aPn2���d����I�͍�Y"�X�X�ޭE!I�=�����>[�\���&@%I��ټ��ԁ�!mj�N�m?c?,D���WԢPWJ~�s��Z���Ʈ@�~�V�а�C������!l�céN�X�{�=e�#���
������������onf_�W�1���o��'W:T�4�*%Ua9K�\7C���)cH�PQ�g��\8	��|�҂���7�U���pr����?����.~3����[4�f�xn�݉j�;��z����j��\�9�;�V<�l����0��>�����N�b�i
�L�����8�`?j�@������?�e���y�(��9Ѵ�6аb��T�ɜ%�'�"�:�c�c]����~6m�
 ���؝��O����M�Y��;�-\M��$�p/>NVe���ܪ���j��B9�_�5.N�󁜝&�Q��-0����l.��KV��ήU�����Nw�;U�Fya���~1�҃u>}ȫ�A��MHQ���P���$ݽv"���IX��z)�.���`L�4b����d�rB��l�4D���]�ȣ�d(����h�CCoo�TI���_u�`nq�Ҁ=kE�1��<S�I爠H�'���i��X�Zз#+��Հg�E����}�!����x�מw&�mפH���d}�v��؍���#�HBo8�¤�`t�����/���"s���к]�E���_{l�а�����v�"�`4�:�a��u�hkEk9'�d/���̖:*k+*݌Z΀�M@�A��*7asK��k��-���2;������U�U��x+E��@����.�\������|�S1�H0K���P�&�!{(�$�9��0/��\+ �J4�!nB�ƅ�%W��ٙ�5��;W�3�D�X�QB���B�*jg�U�������zIsM��*�8p�����ԓxplY�����j���^�����;5b�>��d���h�˰���{̷���J��ю��4��1L���X=_W���h�J�k]��jݜ�Ļ'<��:�Z	/�4�Eq�kF|IMO��W�fO�m� �"JQ?co��(ݰ�Q�x��k/u��p��u Ff�/�#�8�i���ʹ�n@�C�Z�b��7Z}�ȡ���s���F��'��c	�ձI�7����y���R���9ӧ�5^n#�[Jq�W �k�O�)f�Õ���**nI4��(�Y���5��[_�#��$&8h��Oҗ��:Os�Bœ���|�� �`4�i���}!���0�T�3w�K�N�}
�ޮ�h͙�"��F��ò�C�@��ܼp���UH����	�|�B�zl��c��K�zNB�P�/�fI��ɍ;���A�Qf�vt�t�r��Lqi�|�b2�V7�&�^��tC�R��1�V���{�U���:��9�e@��!S��a�8��[!�F�8�"7��wP*�?|7{%��^��5G3��q^�û��f�}���2���*������f���3]�~�#73n#k�a,����%�k4t���<�w'#f���^��?;������)�g�S��y��HU���+M5:c͢�Scf�h���,��`�0��3y�H0���L:�U��M�n���{d�a�6���K���s����F��";U��>��cV�$�`�qM���	��u4I}��B؁�ă�}��Q��3Z]OZ ���s���Mnc=�e{9#����6r�mJ��mo%��?h/�Z@fq?h����[��cH�#FM�X���]$`��R{w��Ny�����)�ӊM��1��i(��ڢ��7�CY��|��C�����Goy	j� ߋR��`Uq<Ld�.����bp'ǃQ@�{`d����s��,����/��S�xG��sJ�c�|\��S9	�O#I�Ea���3���%��	<����J�u��-��cѳ% F����"Giw=ۑ;M����0HNO��b�pY��*��®�%��C�!�
�LЂ���?�n̜�x����6.�~��ՇG}��g��t+�Y�4��,���`����5��aR1��6�k4]�^�)F��U�Q��1�x2���/�K�u�X�ڕ��_���kLDF�!���M�<�l,�;� �nE����#�#�k�<Q�Ų��!����NF
��3�$�
qB�]z���Q��x�N�����}�/>G��@L����Y��c�"<C�`���{��mi���:�Ghz@mT�R9P����Bm|ug	����_�cb{��P��`��BG�fI)m��\�0�R����$��4[J�D'�H��W��1��`9���zz��@�P�b��QL-4�v;�T���x���$p���'`�� ���:J�8��v��g�P3��ƍ ��hj��l���Qr�7��������sI%�N�5�@�0��4�O���R[�?Y�!��e��}z����� .�<"g�ٻ����X�RF���3e�(	sI��l�Uf�ep�g�� щ��-�֠5�q���T'(L[�m�Elyy�.[����M{�ޙP>�����i>G�L���/���N/�P>���|zȽ�=2�6|�@q��7,^v�9��7.���>9�*C{��)i{� �4�i� e���W�\��$��M*�	��G��q�ڗ����i8aX0Z��v'�"��#R����&�U�|���/�;�l���x �R��m��� ���ɑ�Ý�������:AZHTڿ/b6H;�<�R<�8If�u藍$	�[8��d��N��rw[ٜ��B�Ӿ@��Jڝ[y������R;}�B>=,R?�&�-`�_Yq^��f����QH�GH�n�"۟�(���*p[�{́9������ n����' �$�F�Ѫ�W*�Vr��B�&ε{0�$Pd��)ڳnm��a1����%U4�5o������0�R��Uj%9�\@��|"E̚��y����L`\�$�����a�Ȉ�y�;��>�ٲ��Z�٭��j9��#���+`c�5��K���L.�|۾�g)n�i?h�����j���Ԉ�h"��rG(�}Y��K��K�wSk>��K�X�>��C9s]H��d�;]��>�3�N�&ɰ7�h�M�j�8+zW�����˶Z"�"to�l���؊[��;���K����LTah���"�Vh�J
��BQ�ǹ�$U�.X\V\�ry�D�8}�Z$��E���1,�O���{�7I��e�|�eX�zK(J���=YC�J��3��
Tb�6Ҹ�^�QA��ke3u�l�Go7ƿ7:�Ct���y�T3
�ܻ�hR�l�̺F�$�gl�5�7��E҇���6��N@�l�V�"������B\.��?vFNg�m�q	4�솠��j�Њ�~�޴	|_D�5�� !=���yF�A5�p��dT��H��*�
�>֠L#�Kv^#nGϹ� ���ZV��������0�VѮ7 "��">�%��N�R��-�K7���,���p~]��8��^¡���Q�����6� s&P�٬d���|8��J[�:G~�X*f�E��d���!����w����I��2{��&��|����2�����_�$��1�Y8�~@*�gҌ����+��"*5q���<����;�p0M�Fn�51_S`3D�����很\���闚�����ΩW�)^j2F��<Î}~�K<�k�����!�k����61Cr�Οt�'�qY��{�,h�#Ax,0����U���:�݅X+�����:^(�`L��1ƶ� �;��H����܊l^�(�"lo�"��v���������\�o:�6:���,;58�����6�0�SfB���"R��O�8���<��d�.�������X[Ju��9�S�r����H���H1޾�A^�"7g��x?�I�� i<(�؂��m�eօm�}Wi�� ��+�L��R�������k��t+Q�/�xD�?uD~C�K�^�$v���:^s�t�G� JV��`*�5�'�D��R��]�Ƿ4Y&˴����ZÜ�cZ����r��tr��0��{J�j�s//:� �r��!�f3��:EkA��������]���d�F'�,��)�2d:�%��6gLC�u6��Ң},�y���Ј�NeFFE�.c�=c=r�n�\�IM\|=_�S�Acy��^��m&���GFC�<2�Mٙ�E�5�p�o�1�����L���v��3���&%	�7yM�Q��%V<U��99�#�\�� j@��z����2elOO�)j�ܛ�x;Y�$�p���Ub��y�fβ����¸ݵ�1w�HɁ�G����&�[��k����zWߛ�5�oQ2_����6��\����/�$���5�h�7_$"1���܇�^�9oe��7Jd\�p�E.�iT�L�{v	7�5s�rk�3���J���C5�@ȁҍ@o���?��8Cz���˗i�a�ݝ��Y��d�m��X�dtu�	���0�BM�k~�G7�'%e���&.��Ӫ@�]3��gʎ��_+ѩ^����c8�2����HFH��d{ �5�B�����ڮP�K�B�	H����|�T�r��8ؐ8���۾�A���(JfE���8P{��("�}�V��d��b�g_f_�p	u�̻;^�9�D��0�)���Tϖ�4XO P�m�{f�*�9���;kg}�Azq�S�l�WO�m�����*e#$��x��`���=�E4=I�j?^�-'G��{e�bM@o@��G�&���b'�y��5�ģv�;u��L�ʥ�xY�r��H<7�d���悖b��B�w�R�*\�'\c\�L!���A��˵ȅ��$`ՓA��X�o�����������Ia)�!%��(v�����C@�W5�NQ֮���C�r׵ܝ0��d<S	?3	��L�Oၭ%ې�C�]�t�9f��(�e���C�i�m���M�
�Mc�+SśL3��5p'K�/-mt�������`4��3�
A
�1Pa���i�����=�%��Bþ��4V^;=�g���m���%%��0lW7`!A|8����#�n^F�>-	��fį�v��6��|���2����p��V�66�Dgz�׮��3�>�䨸�>�V�b�����P��84�5�F�h੝�K1�I���<����Y���n�P�B����Az�O�����N8/߂�+�CH��MZ���F����u��~Sd�m���������zd]�q9~At)�6���?ߑDK݂�Ԉtw���e5ٸ����djvç���b���2op��-���YUC���#�A2�}x	/tڠ�	L-Y��%L�B@��"���r]�Ox?O?��	fB�*�R�0�������aqxnޤ�?�y��Smd���wʈ�#R���kmn|F��/�}��N�y�U�k$�����;�O��O
G����DWx?�W��<�tfؾخ��VT�k﮴>9���?�U&Y��w$.d�6}W�?P�rP�ݪ�#{�+��3��x!��R�q�X���"|�-05
�?y��z�(�h�V1��� P?�B�S��;;!Lţ��a������I�u>%p� �>u��Ĺ_������a�y51�{�^��=/h>-D��9�Chz�[���W�H�}>p{M��!5���M<ҤMӰ�U)�l�Ը��f�O'�:��s �����R��bOCZrWg/3S�˧+pKwٿ�2�?���:��ܐ�eO��&�ܬ���RX�Q&fZa�<R�?ָt���$��̱�
5!�'�ğAɟf�j�B��r�mc
<�'�<n��q�0X�w���(0�%Ƽӱ�PDי�H����=��j��f�H�얶e.������H}�e�Y�!U�M>`J��� �Y�@����4� X�E�_�E��L�W�U�emIϡe6*��諨.���Y˥�rf���,���S�����4y3��_���l2���z.��P��Ƈ|+2Q`$��Ԥ���
U|�T[eKbɠ���TI@"���p��&�Y�(1TZ��$�#��4�Q{�̰�P���_R��r��jI<Ќ5vW���ޙ8Q���}�MW��m�ޫ�3�ad�7XnB���t��i�b�ƧǊ�BEBL|�B���A��wyV�b����	dK^�þ\�N	<�hL�鋆�h945�D����u=���'@�ǥ�o���ƙ�\�oe��� ���Ӂ�V�4Y9�/;��ҙC��`�g2&���H��R�������0���a;&�m?��.jO�@��FQ�;��*�G��C��,����#�u���<������X�r�M[1�*�O�50@�4!_x㶱�v*��Ug{��T�ϋSl�~�dIb�jx�M�t�Q^�p�"��&ߊ!�1�ӫ֑t��u�'i���۱�)}�7-u��9[��UZ5�y-���+�����%�#c�=�I-��\���ͱ�zCRL�=��}ߏ5�R�q�\vT�V2�-��N݀�xҿ��T��&�Ϸ����FJv��;�g��<�VO1����8FqF��d�������f4)�x,0��H��Ub�u���ګLW��1S33��1�tS	�(��!����\�eBOl�:�of�7O},����(������$J8�����$����z(3�"t��h�����8&���4���~�÷�t�\�'c7����c�ZV_`7�xF�Q�K��B`D.8X�%5�	�I8����DO4�OD˪��,}���������b#�����wr���z�5qm�AwGzP]}H`���|��v�9�4�⥡'Pk�#WA;�`��g.l�
���@9Z���Y=<r@�I���ݲ7�CSay���Z �������β�/�#ݍ�$�����'�ͩ�Y�/����5����	�V\��1H�3�f����	7���}���ȣ�h���y�v�s�a������D`Qx73爏}����Ny��b�E�@�X`�(���ޱ����qn���D�}�#� .폊�j��$���.�������?鷆�#0٩|x���a�L���(_qǧ�`Qz�d-�>!<G����v��zu�1]�Mb����߅U?��%�[7�?���eT/��V�[�}ef_z�g0ݐ�;�b�ݚ�#4��t
�7���$�=<�(V�^��f!�%�r+�u3(��D���J]Q2=��b[uC�@ή�	��jW�g�h�WQ��+�$�����g�g��6fKH��@8�,��G����>~�y"P�������$�XL@۷��aO�f�ߋ����l~eζ_[
�j�:�fG�UA%UTȌ1�6lb)莑����������f=�ne���~�/�R����6�?���	���~�!�b)�	���֩G2f̿r�26�ĘP��R>6-V�Z�����]��8ÜS"@ۍ���ݥR�|�R��b�F�pn�{lw�ڑ���7'����#�F�D��h=ً��
(�%0�B2؉Av!����eh�Ǝ��=��>A�[��h� ���L�X@Jn]�('z��`�q$2\�iMx\X� �2���d�F5]������Uy�*�=	5]�J0�^��j�U�I�R�JY�8���� х���^�5,�gLI��S�|��F#��N����u"/l<�&��9��S��8&"+���ͮi�t�ѭ���e4���l��H�2��+�E�).D	�Pnu���f���^%B"־����ck�>�����@�6���P�#�������p�W�ne������n�H���9G:l6��Ʈ1�u�*�;�{�4�c��2/�*���u�9�P��n�r�dC�$�ケ�6�F�Prh�l�<��\�FWI~�aD(|�&��j��
�4�%r�8j&�;`�l29��D;%8u�p� �^�������������-̍j}n����61����G��R��#f��p�4R�`����
'��.�+4ã^���� ����I{��yDv�\K�K啐A������Vԍ���0�S���X��dB�z��쌼 ���*�Q��c��*R�2��6��]�|2�DG�`�������⃉`4lHrk	�h��|"`��m���i�3� ��R�\�A	� 8��^~��L���l�[3��ǂG���Ʈ돆MP��j^�"�<Za��h����~ՙ�C��D:R�ġr�' *<j@-�;7��%D��y/��WO�[������(ʡ㛵L�u��^=�:�*�^:a|�S�#�����39�;]?L��g��@�y����B��㧓���%?���7_�%uō��\V�{K62�	�.��#�]H3J��E��hH;t{P%��=1B'�1�D|%�W: �0��㢯 z����@�Ϙ�����.�i�	��Hv��>3`�raM�;��pS�?)�~���L�E����cX"�v*}/n��&�o
b��qZu��8�E��,�n�O��}5.|"���s�3��$�,�堽�j ��F�����D!�٭�_�>�%�(����ǡ�$�jE}�r�܂�,�l�[P����;f�}h�ѿ#X�E\i�Y���c�u�n�ь�u�{�[�ÏMc>�pB���w_p59��馹���L�v.���5�"�nF� sQG�g|$����`vu浖��G�m�`$A��r��������<��L�\�q�9s>�C-&?bA;~m:Rg��A`�/l��ww.���9����w �H����DK̛IJqx�!�M�R�s)c5�^�.�q�2$��שԈ��g�x��ω���|�7�A�YV�:�	���e��;2��ޠ��g�:#��m��<\�-��iETN
�o��a�2؂KM���TX	�����:p��S�k���F����Ч��N�Є�Db̸���6b̀#�������syЈ��7WE%�}�����FY��ȄT�oD��;O�ǒ��9��@��������ve������~u�F}��[�B�@�|�_�;9rH���
� ��=��]�"{�၉��_�6�^Ў���X�P^h�\����$i!�c��Sd�޹'�z@�]��J�bk���n�5�ٺ���2C�[θ37<�P?�0�Bo!E��rL�A��hwgHm���c:T�癣��4od줿�y�F�
O~�:>�I	�x�{�4��E!�\��_��cu�C!]�3��T�	Y!��T��X+r���ǴK����%��������M��!N��B�p�Qʫ�������K�� ����m�z-W����kF@Wt�S[-��IAt�b�6�{�e��n�[ye|�um�����^�{KA����(��o�=��4��e\mB(�RF�K�Y諟UDN��t#�`��]޹
R�O�hHR
�����*�2a+�t��C�RP��U>���u�8F,8��`C��MX3<\�-��e� "�V6��������8�7Ջ��}���O�s���Nؤ}.�;y{1Ll������Y#���;�	`b�Ӧ5w!���瑯ݔ���H|�GҤ1qNc7m\�;�2�s6�$����axivI�r��mAr$�����5G1K�:	+T�;eՙ�ե�w��&i���@c��s�M��� ����ǜ0גTь�]^ki◷�"?pR�Y�p=�5\V�J޷�#*�r|֟�?%�M'L���=%@֘�3���	�����9kf.�-Y��vk��S�_	o�{�;����,K��Xκ+l�z?p\��$>`$�s��I��5x�.��B嵚�J�3H�{�T�$�ؤX:�6�&�� КO���G��r�Ǉyk�� K��4�`�>ű.��	��,�?']��;hg �n �Ч�
�Z�X(� �����:�,�&'^2PUӥ��)�E[��WM��ރlNE�L7Kԫ�in��:i��믕�wZ\�����ű̯����Ă���j�]�����C�h@Z��^ �@���;Y˿�.��_��3��?�з%�̻�r�3��ڴ�ŏ4��������ٹ�i�}�7�1y 9�c�RT��c(竱� �ۍ�?�IL_��5H袿�A8���P'��-O�&����4�ٟs��Z��U���w���U���G�����ZWm��O���V������5>�����޴Ѽ+F�F���6�湋������@�G���ԋ�cs��ԟu��c$��C�O�0�i�ƅ��Y|'������_���KkM��uX�X@�*�-��Ǳ�}eo���1�4���a�e-�^9J=����[+k�]V�\��žo�i+�ڬ��W2��^�j4�df࿷�<<���kj�;٩�(Bqp։j�_5I�J��Z���N^:B���c��P�CC��7#��$$�T�7�V�ӺO�Y~�q|�fS��@�k�;�FDѨ��ң��^M�~7���'�C�T a�����r�8>%�}����p���>����͙?S?� eǓTT��f�ar2*=�!�����g?������N%`��]tb���n����R�8�֦�K�X.q?�B;����c4P��?^Q%t�a���L�D��Q/��K�So���%<۔%�B�V��Ɛ���n��f��A�B$��ǧo7���b��T�n:����GLi[_�ܥ{�f�c�[�kejW?���f����uW{_�i�'�`,~&�� ���u�	�qe��Z���I[�ۂ�)� �,�c�F������Ei�����}C��F��lN߱���i���'�ό�Aw2;^�a^�=�`u�%��r��C�`S���s>6]�r�Xڪ��	-������CY��օp�.P3ٴ ��MeY�j��A���}��m�kU�qt_�m�	��抅0�n=�%�2jHy_����}��vۄ�x��UVqc����g:=����Y��y�B��x�,V�2��n���I�#��͠��$N=�.k@m�ڤ�}�NCY��i+��%��F�ձi����G&d,�S :�t����!+��/��@Y������򻧲��kp~�:m������HiJH��&��Cl ��4}EY�
է����bv�w��p/L\_��q����#�ζ"S�^�#������HLQ�L��{��y�q}�${@R���k�8�&��OYg�7���T���z����t?1n
�X���>W�
$4om�r�����"�W�i��p}"��g��;�ڝ�DO��i�[x�,��UuUL.��?4�������e����h#��8�9D���4���o�`�+���g�gh3oycUA�y��G���l&^�[Q��-�T�L��iv[#N:�	�d1����.�oT��(~S�ͽ���S��$��v\��bw�'��fmX�bߨ���R/��ͷ�c��N�ٷ�w����x��ee��	����۟޺|@w���	���ji�mayϹC$�_q��k�������w7}b��^�����Y��%��u�ٳ��ڢ�M,bN�~� f��F�]>�d��'����յ���˵G��n�r���L���P��ZR^]Q�c��ڭ�Gl��l��Sid��H��:��Y���+�&|_�[LO22xĄJ�:��lZ'������c���,�f!�S�Es�l^@K�����Ϻ�q|��'��⊧x��8�||�v��5����ŷwZ�a1[ЅKϫp��I���,t����ڴ�ݯ�m���~���:�q{c������Y0��1��C����0�.��t�;��@���x���:�7v��$+heʅ9���Sn;�A,�5vI~Dς�N���ķ!Q*)�4�I�T�6�L�����X�5��M�֐FóJ=��d eU:�G�?�K��8k��9ݗ���8�M��9�0�?�g�>�
��x5�f�5,�fs�`(sX�I	'�[�4��~�G��h|ik�8��*�d�]"Z���EE
c��K��o����+��O�5�	p�Z��*m�7h�<��c��7���:K3UH�>�I�>:�=A����kgɦ ����u~�1����{��xn0��yW��PْR����|X�$��A Xh �p#<F��8�b�P���^}ǐ2k���	Ҹ�$�3�,
�C	黟5�,�Op"K���➭�wG��7��r��K/>Jx��vF��v��vGW��
��2LF�}�=v�=���B5I.����[D�8�e7�OnJ0l͂q��a\�=�Rбٻ�Z�� �.P�#�����#jH���XK*�z
��z��$�X��x��]�a��%�w7���)�\��Hw� ��`>���Z��˃����
�}�r|\��D���֘eL|h�XFrȈ��K\��y���ös�(��LF�#'?d0�������w%d����{L]]A�
���GO���ƱF�ei���s�Lv��5���R 1�X�Gw;O������t�՚D�3~2(�n����y���
*����g���[M"^-LԖZ���\\�����x��Pi�=2�q��2!��0e�M�g!j_��XT��(G:Ѐ��M���L����R��l�K2�����K��2sf�Yf�����X߄��,U�4�V�zO>n&�v���Ț	�����w���u�>�߳�?�Q�T���Ejn��-'b�*ͽU�I��~��PFf�0*tx �/�cP�'q}zM.m;Ew�Kt%*H�7����o[�����*�zp�R���O�'x�Y�:-Ř�;��x����]V��vP�1غkDrq=p6�y��N5b�+N���[9���� �}���!�%U���I&�����_A؝f��RMs~�;���_9������}�H����O6y�|�L�O�:����kVP�i6F�� �����x��jP�m4�lV"����bۉ��}W�>uEj$v��S��T���,���T����E굋 f�(���|�-����(��:�#�=\�m�Q>�� �]m}�? �c%3a���9��9CP��_z��L��P[�����Y��8�b00�,~h��s��T�p���B�DT��#�3�L�y�
������C�Κ��M�����"��O����Zj���2,v�3�Y�v,S
�(t��XsX랚�z����+�:�"�9|�6.��A�$���=��U�d®!����; ���G#�Q��}�<���m4EQ��R<,UG�Ti�S������U�Q���b!Fa��l��_/�P�#�;~r�R��XP�� ����GB5��l�հ3�u�S܀���D��1��6A=2?�����R%��Z�!ʆ�-E��ߑ'Ӏ�jGn��H�WxD�dA�i�m\詄�+�ޤ��;�C�)��gI��� O��Ye<� �k+��VU�,�$W`7��'�(D�4�2�Xb�JJO�����۪Q�o������)0%�8�0|��/C�ɋ��Nbm��f9sƤ��@�߁.�aG�]��e�t�(1�h�[�Q_@�X�4�ҬN)��-I�4엣/z㑺�Nm��=m_�\�Qk1L<��!�u�-�E�.̂X��
[�I�*���wRA}1�I��U�Y���D����9'��h.��7E�!`���d����#ky�W�J�B����2'��Y��A���P#�=�J[G_udhOS�`��Ks����Z��&)����B����5S���	�F�� !߿���_Q,��&�w�]%{�x�Yթ�5�2�Ĭ�ս�H�{�\�?a0�G��=n���V��"�*�����Ȧܩ���Tl���Հ��6�,������y�{�`3�R�)3�h3���	s�`��tU���-X��VŞ��Ơ���h��nq��'��U7�T�Y�%T���ݳ�� D� ����s��R���4HE�)��k�� 	�q)<XM����Ē���Ybֱ2#s3xs��P�Ox�Ҋ+Jڤ���b���:��HOKE8ِ�z�*ÃO�$kar��a9�'�y��Z���#;.>�7&v�_���iΛ7P'C���+	=��������Hv�R�[��j�U��N{q{�����̨\�C�%Du��c;k�KXG?��ԓ6���媜�?���#�[O.Z�pQ��<sf����z�>WG�/�aP��,s��:��$lnKMĚ������j�s��I������u�q
��JaŔ���ƃ���B���-���4f��)� &I���6!,7x2)b(�нu*R��@`z�89�~l�v�J�f]� �����Rx�?n� �d�Md�~�����\%�%�Tc�zdp�@���\�Q/��a�V��|�ł%��[��ě��6d$/-o�;Y�4��B�G�׳[��d�e��Qf�xY��Փ� �Caԟ�O[,��v����2��䁩=��)�#�l�C�-�]�h6� �ۭ]�����~9H��4?���~���p�6F��T����#9��N�ʨJ).����}a6K�綬Y�0e�~䀶yː�،8�"3�M��~�^��ѩY��.F"є��8
�p�f�>57�������j �(��A�m����	����:�E�&�o�p%��	M�X�:�n}[�d!�8���"�ߚl�Զ���(w=�������}P>D���T@�*�Ma#�*��x,�m{S^z:os��M[�MА�� m�<uJOL�v�����4M`ռ�xy�K5��?h̜�R�n��U�㞟=ㇻ�Ywn�������=��x��Y��j�̧��B���#�fL!����!ߨ��E�ze�%��,F��y}MT��U�zT�����b�w��ee{��7F{�'.e��aD���ǖ��y���ǥ����~(Hd��?L�(T�o3�1�����WT��߹z*GUF��y�[��7���٣_[���y��0�¾�\b<��� �y�?�&�">���	��d��B�CM>\0|�o%[��G���°��"'�ie̤���B����g��%)�%h��I��.�V�����HA��s���l�b	�A�Xm]�}ٻ�,.���V���J��lv�I�*J�W���6��#%��N�yR�r��3`7C�|�\�p���Α7�,���PG��~*��/b��MG�,x��NvO�+挤�Ό�Zr*	��xnA��h�Ku�������r�g�F	��6�cdn�a^M/J�Ï������3%�pm�1��~�#��s/��6ڄ����;(�������5Q�J���Ay�F�eL���+��4~0�ڴЁ;'�{H&�V���	"�oq�V�W�s�n9�|&���Ň�6���u�P�rH�T�9�ɰ5mve
Yk���E�X{��~�$�v�C'Q�W���&��ôBkX����/��<���.d۷�]v��u���=�>��I!O|%c�u�M��ѫT�<N�<�;@�$�)��%t�y�LD1g�S�a��Sp���k�eZ�b�aFzR\�c.�T�o��v��|p��!�>S���+�0��aPȻ0��|p��	N�����lm�D�貈�ʘ���P�J��X��` M�a���X/fmnw���	|�a1��J9YQn�	�	�'T��~0�������h&�dXK���Б�y�3�Н�%�:CC:�>"i��S�P��يnF-,g��*�RX�;#�o~L_Nq��2��ma:�s�5�{�H�M�Y	�q~LE���X���=�!���d|� 0�x��hΦҼ3'bfT@��!���v[o���JI$������Wʥ��(��;��;,-�6������|�|WC����럣��b�����;hqB��1#��.	_UO.�5�`��ⶥ[bc�%��M�ĭ�R�Ĩ��
ǰ�r�3v	����F����^��(
w�m�ׁ�_����pD$W�y�O�	�<wZkOQ#��j�?LAu����",��8�n�+����.c�'c Nc���H�3Yw�I�����ٻ��)	D���w����ڛɱhYk�?dDf��aI_�\��[Qw�$�jwUd8��<�����6����꿰V7��κ��b�4
My��o�n�f�c��� �Zk�����+H�E�.���F��ǶM3��]��cv�x�f�|���������[�9�"E��Xs��	�X`�K�Ð��Ԣt6�����5,5��$�ƭղ}58DC��d�H��GΠ�ֶ!kp)d9�<W�\;����*#��*��e�Y����K+?7�rJ"8J�l�L�v�u�q-���1LV���YU�W�Ij�i��|,�?bx)�>�-\}�^4/<�Y;�֤�����de&ޖ��g���gN���P�p��q�ȧ�(�w��9�c_�������%�=���҅�J�7a����M!Z�/�����buE�*��r�ME�񏗚��^6��0O�Piu+v���z��m޻/���qi�|D��h�ѓ����{;h?�	�f��Ӆ"&�P`��`	X����P��Co���Dɫ��"O����e#�	�æ�`����������^:o땓ݙCj���>��4S$T��3T[�'V������H#�%�ZwG-T�-JS�m�ƪ��>ۜ��or��^��c�K9ވv������n�9��< 6�E��hL�w��e���-����F^>��o=��j��TJ�(�r����41C��Qˤ���l�� ��R��ib?\��풝]��0p\C��E�u� ���n?��5!��g��H�ω3yv��&�SIO����B�͔��A��uZ�%�i�<P2��p	}�d|���Ӯ<t����is�veX���Gל�$8��vh��$��P�[�[B��.�ReV�\O>{��T����X�F)Xr��H|_�.A��w2��Sgsg������Zs���F0|+p"�U���4ő�A���}�K���?�C��;�M�)`��1.�j�j@["3���:>��x`�E3�}�s��nuU�Dp����p��t�(,�l5��y�4F�,t�E%[0f�@�}m�sc�~\��8���z�4n7�\��2�(\3�Ծ�|C�5�\��\Bf�VK�H�f<������D'M$�����pv��+�\��7�cj�M����\�u��/��
(��Y��\��O���8
u�dI�׺ݼb�����II��F��Uc�U��C�4�[����8su�x{���i��M?>� 7����jb4΁}��:�3 ��bn�sM�@��%k>��T��@8\zH�ɝռ�Z� ����_�#t�B�{.o���{ޭ�%��L�P#G�>��ϫ�3.�fS�^zm�����Dy�z���E��p��!���9�����3��y6k{��eA!&�^��S;�r��r���p�3�+̵�tJ()��d�~Ӷ)FBS�x��cw�O��:��Yy��w!��d�����^=���)��Nֳ�_�H~��m_a��QhI��Bͥc(Ѹ���u���0���#ir�T��ˉ�����k��v�LN� �>�|�J���!I�PM���Al
~+!s8�C��xh%�e�(�X]�Q� p_-�I\����,�,��d�J��rSl������;��`�|^��s��Z:�a���Fn��������^���{.���K�k�W��lD����~C��q����+����_��D=��/��"�����Eb�#�����>�'���>��;�cNع���e�ÿ����Ν�T��9���%�X:�^�S��N�{�@�ס�F��/�;��>6���GMכ�쩏zS=�U(��>�|-'�uK8hFW�iu��nk��g9�|�N!b$�����ѡ-��������>�@FHB�gQ���L�׼�5�$k%b54���z��2 		d�E�yD���K˥Q���6nĽ�Xu��2�=�j�<T�tJC]���VJ�|~"��O7��ۻi��A}�V��9�Q�D��ΞL�t&�M/���c0���Bh��DҔ3��fi�k#(��H������8�#�"W6����!bR�r����@��e������I�`����7v\������L	)�%է8g�r�*z�}y3��������Ϊ���URz�_d��뷧^���^���a{�����8B��hK�l�}S��뎙�����E�M[�^�$b��:��؃��t��	F�NXk��XP��J�G ߜ��g�T<��Ū���d���S�:aʜ�al��Q�Lz�xv�O�Ïov���p֗l���޲p��$fو/0�:�TY[�	��+j�c�#�n��3g�ir%�j���c69��4Y{1e�_@g5{������1�Q�]SG�B@]��JN��1Q�f#��΢��vk��� N�X�V���P����K�.�7���u�� �=b���,��wi7?W9��pܣ��[ISw[]󆷅`���x�&�-�E(h�@`l�H���K�Q���@��9]l5� �T�a#[M�ѕ}B���t��:
��>ס�fVA�Tǭ�B8��U��sb�p6��>v��i���D��+�Z_ ���/&&��@)2���:�M�O�+��*h�-pn�45f;�C��/:rg�����q3��a��b0�ߘ�2g�������l���A�(Z�a��kA�ꁜ5ߺ��"X�{f���n�����u�m:#�p������^j`7�g��Hk���zz���J+U��B��4��sȞ��^�%q@��s}z��;�rE�,�6�qig>:�n'I����-V�rǾ���6���2=��k��Ls�\��ƛ`��O�vJB$,8���j�1�B*���d������-���������d��bR ގX�TnZ���L�۬t�#�)������X�S�Cv���icg�fO����nB�T��sȐ����1��T*S{�S�3�.��t�B6o��.a��g+~7�o�a�w���x�R\��pa�&�I:$@ �<ca�~�D��[L�+D'Ϊϴ��Ϗn�=-N�"��w#$ʪI}�7۟A�YY6�_��D�M~qg�O�p9�Kp�1� ?��̡��`��BM�\�Q�>��2�����/C��3S.�	vhH�U
*��'4�ˍ̣�HwP�P~��M��3��1��cV<;��u��F�L�ꪖU�Wc�\�r981ku������) "K�H������oZ��� <�X�W�O�X�U BB�s�"�� ��9U_5-��-���Jxo��H�cr�P[����(X��mM��9���T7��\��ƜȆ���8!���ΐq1*�2j�	z����G9 �G.���m������%;N�.�Pщ`zfC���Y+�I� �#�D�y\�#��w������x������רw���x����f�\Rt+�K�;�E.���}P�!妋�Z��N�e���TX\x����s�������D<Y����J��q����I�${���+nQ7H�p��7� Ͽ�~����7ט��l�8��"�/��_�x�dr�}�=����"Pf8'�Y�2��^�U&�'a/�,d��Q����,s�\G�MGF
}�D�Zَrn�h�}1����^w�<#�|���H}��>�ps����s. e�pW\Bz� �>�t�ⵎB*��:nz�������=i�tǒ��~4/w�j/
� ��������1�����ah�T)��B�H�v����y��pۘԋß�'���k�B�]0����rO����֊��5l۴š�$����YSz}~N[pr+R@S�1IWOɱ��@5l����-ITr��L{�G3�����cg�ZN���6��/Vu5r���֋��J�޻�a� ���u�y;[�@���@�s�>6J�D5uH��O���E��28~|�z�E�H��#�zV��>K;���rxj��k0\����:����w�L�&�J0���D�TI[�!��j�ki��j�`�z���g�<�WW����m�:í;�ȹl/�.�!3��Ug#�Y��i���[�C�6��Q�dm~D��7|$�Z2�����Ж���.��:^1jIe�Z2���8~�y
w|WA~��Z�q~��Z��!_����������:�Z�P�᠓��Z����-������jm��hW6k���Ũ�t����H����[`��|�?�:�z�A�|��Ki�W�̡7�M�>D���jѓ�p*uK��mq.�3w�C�@� �Q��t�=8�ौP��ڟa�e)����~��.������R�����{�ѷ��1/��R���4s�����k���7����Gr�P�2i.�<��Q8J��=�̝��0�_�Y�|����;,c����Y�7Z�Ry�1!�Ĭ��� >�'و�>CD�.N�MT*.9I��륓�
�&a>����桼��JW��(���])����4��ۖ���h[.�iR`n �p!��uV�2�:�d����Ա��;�巋��쨛o��XIr�V�]���&C\������Z�G��@��<�9 ����P��|�}5ݎ�i�c���K�EKڥ����8/&@9EN���Վ�2�����#z��b� #
���,������%���ض�;v�|f�ʺ/|�W	���S���Ա}2O�g��b*;�F3�%6��F=�s$���[�7�����8��[��?)ɍ��a��*e����f����Y�_��Z3l���fh��?	T�����?ߍ�(N�b�4���{h&tm�6_�B��pqY��*�8���:nF��#��h�kos&~F����]$|�&�i�X;Pq$ݔVӉW`��LJb �b
gzځ�Z��K�����2ɭ4�g��2�ñ���{I�'N#����{*�I�k�ݣb��r��>>]1�O��@V�$���QBɴ��:�5$[��ӊ<��>��K-�4k0�q�Rck'���o������\�H�s����D'S�g�~���2h_n���V��@K3)�N{΋ �Ю/���x@���p�_Yp���T��Т���]�k��ݝe�LX�ً�:Oo}� B����B�5ǜ��aׂs�N�C�����By��v���V��-!gL�-0� �A���� ��	!�W�l������W��8m�U���W���Q��HA�!��D����k|rQ�4^f�GP�+-��1{�!�j������d�	*��K^���8�-�*ΐW!l�q�*��k�v]�ZӼ����X�Om��"x1�v(츀���.�Q��r� "��zO@r�{k�vSZM�A��x�
�Y���P��N� ۠)5��xo�4?D@ͪ���pS����S/��KpN�0�+�k��S��=�P�s!<��,=��lm7�:��?<Wϖ9�zFAVy��H��[v�(�z"���e���_>ب4*1YOk?Yu��묦tm��ȋ�Zm�l���#	FLl�4w�+L�t͌U{r��Lmz��H�
#2�"��T0ҿ'�ndCsV`��[�0H�$��m��=�q�Ex����,(�{`��'���6=ʮd�@R�刵Plm�^�w���/�<}�zŜ���x���� 19�|L�Q9�����im7V���S��r ]H��4����y��������J��
)lp�$��Y�Fw��+��VT�3�=���8쯈j�f쭐a՛&�f���,��^�o�?��WW�z8���7���n}?xǨ�%ԣ&�2��І�t5W�߳��ڱ>zʻ���k�7�.�v]7���$�*O�7���zi��:	�Ǽ��&y	Y��e��tJz�5n��7T1�=��ÝS�as�ͩX]��tsP�R����%�k�cF.���6li�t�y+]�56�,T�{�3���؊��@y�s[�ڂĖ��d�:&ҿ��GN����J	�bd�U�oct$��H<��c�T��oꁐ�y�V����Չ������-�V�nm�]���>3��ikTscF���K�b.�kߵ�\�b��S��0l�̎�@�Pz�Mo������Da�����2��
�=�=Ґ�$!*�H�9���ÃX⣳��[N�<Ku�j{��x.<�Q|t�8I���$�#0�+�s
�0Y~z�=�p��V6��x�7� Q�J-d�\�Mp�I>L+i`/�/d]U��1�ڦ�@�����M,S��[C$ȬٚDC� �-�h�����fפܔ@�l[�����[��R��fЊd��ss{�s�UF�ʥ;og3�F�� �1��s1��2�v��0�V*�,ۻO�gm����+�����|�٨%	t�6�q����|m�K�{����Q���mw̦��Jx*����$�@>��z�K��$<[r����W���=���߁@[���H��Y <A��^��������K��-Ř���.
y��d{XPK��J`���u��5��7-"̞�j��>�i�	m,��3�,�䀯�/7���E�^�v"�i��/�ݼ}�r���!��|b�G�{F�y�l/]��[
���ޔ`>L<�2��T�+9�3B(A�8D��j��6����!��m�e�)�"�Z}����$�"���=�����k�d��فƋF�ߓ:��[�|��dC+1�;�UǀO��S������x�_xt@��pi��|�@�o��\I����B�&M����w	��)XD/���� ��
%i��]w���~�WL,������ٚ�Z�4�1�`�	�aS��<���8��UH�v�a	G�}���e�ڒ�	��_d@i���M.��\# 4RoDP������Ƴ}�э\���R6k*c Y��N����3�'�{�'�a��^�t��-�:Cz"�Z�ʧ��?�7_	�\1(޴�J���V0���S�{P�vɲ4i�;�9T./��V�~�H)�W���6c��k��D��'����B`H4#�^���i,��E�%�m���S���f���*L�A�T5�P��<�;n�%,l6f�XdI̞~��ʊ+���]�*t�H�$C�H�<�QTk#WDa���S�ÿC3��x��6��7򥓌8f